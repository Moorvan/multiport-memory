module Memory(
  input        clock,
  input  [9:0] io_rdAddr,
  output [7:0] io_rdData,
  input        io_wrEna,
  input  [7:0] io_wrData,
  input  [9:0] io_wrAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:1023]; // @[Memory.scala 16:24]
  wire [7:0] mem_io_rdData_MPORT_data; // @[Memory.scala 16:24]
  wire [9:0] mem_io_rdData_MPORT_addr; // @[Memory.scala 16:24]
  wire [7:0] mem_MPORT_data; // @[Memory.scala 16:24]
  wire [9:0] mem_MPORT_addr; // @[Memory.scala 16:24]
  wire  mem_MPORT_mask; // @[Memory.scala 16:24]
  wire  mem_MPORT_en; // @[Memory.scala 16:24]
  reg [9:0] mem_io_rdData_MPORT_addr_pipe_0;
  assign mem_io_rdData_MPORT_addr = mem_io_rdData_MPORT_addr_pipe_0;
  assign mem_io_rdData_MPORT_data = mem[mem_io_rdData_MPORT_addr]; // @[Memory.scala 16:24]
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = mem_io_rdData_MPORT_data; // @[Memory.scala 26:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 16:24]
    end
    mem_io_rdData_MPORT_addr_pipe_0 <= io_rdAddr;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_rdData_MPORT_addr_pipe_0 = _RAND_1[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LiveValueTable(
  input        clock,
  input        reset,
  input  [9:0] io_wrAddr_0,
  input  [9:0] io_wrAddr_1,
  input        io_wrEna_0,
  input        io_wrEna_1,
  input  [9:0] io_rdAddr_0,
  input  [9:0] io_rdAddr_1,
  output [1:0] io_rdIdx_0,
  output [1:0] io_rdIdx_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] lvtReg_0; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_2; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_3; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_4; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_5; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_6; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_7; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_8; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_9; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_10; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_11; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_12; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_13; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_14; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_15; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_16; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_17; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_18; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_19; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_20; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_21; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_22; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_23; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_24; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_25; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_26; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_27; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_28; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_29; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_30; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_31; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_32; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_33; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_34; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_35; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_36; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_37; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_38; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_39; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_40; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_41; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_42; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_43; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_44; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_45; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_46; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_47; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_48; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_49; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_50; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_51; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_52; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_53; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_54; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_55; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_56; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_57; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_58; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_59; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_60; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_61; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_62; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_63; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_64; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_65; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_66; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_67; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_68; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_69; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_70; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_71; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_72; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_73; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_74; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_75; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_76; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_77; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_78; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_79; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_80; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_81; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_82; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_83; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_84; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_85; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_86; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_87; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_88; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_89; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_90; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_91; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_92; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_93; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_94; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_95; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_96; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_97; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_98; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_99; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_100; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_101; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_102; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_103; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_104; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_105; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_106; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_107; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_108; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_109; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_110; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_111; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_112; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_113; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_114; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_115; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_116; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_117; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_118; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_119; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_120; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_121; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_122; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_123; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_124; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_125; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_126; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_127; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_128; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_129; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_130; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_131; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_132; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_133; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_134; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_135; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_136; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_137; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_138; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_139; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_140; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_141; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_142; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_143; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_144; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_145; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_146; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_147; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_148; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_149; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_150; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_151; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_152; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_153; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_154; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_155; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_156; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_157; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_158; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_159; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_160; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_161; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_162; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_163; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_164; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_165; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_166; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_167; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_168; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_169; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_170; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_171; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_172; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_173; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_174; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_175; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_176; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_177; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_178; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_179; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_180; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_181; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_182; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_183; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_184; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_185; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_186; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_187; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_188; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_189; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_190; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_191; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_192; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_193; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_194; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_195; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_196; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_197; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_198; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_199; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_200; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_201; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_202; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_203; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_204; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_205; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_206; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_207; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_208; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_209; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_210; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_211; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_212; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_213; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_214; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_215; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_216; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_217; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_218; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_219; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_220; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_221; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_222; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_223; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_224; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_225; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_226; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_227; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_228; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_229; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_230; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_231; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_232; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_233; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_234; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_235; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_236; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_237; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_238; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_239; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_240; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_241; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_242; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_243; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_244; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_245; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_246; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_247; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_248; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_249; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_250; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_251; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_252; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_253; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_254; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_255; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_256; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_257; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_258; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_259; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_260; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_261; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_262; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_263; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_264; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_265; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_266; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_267; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_268; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_269; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_270; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_271; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_272; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_273; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_274; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_275; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_276; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_277; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_278; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_279; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_280; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_281; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_282; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_283; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_284; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_285; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_286; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_287; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_288; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_289; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_290; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_291; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_292; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_293; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_294; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_295; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_296; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_297; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_298; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_299; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_300; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_301; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_302; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_303; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_304; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_305; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_306; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_307; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_308; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_309; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_310; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_311; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_312; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_313; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_314; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_315; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_316; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_317; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_318; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_319; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_320; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_321; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_322; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_323; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_324; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_325; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_326; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_327; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_328; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_329; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_330; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_331; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_332; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_333; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_334; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_335; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_336; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_337; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_338; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_339; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_340; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_341; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_342; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_343; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_344; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_345; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_346; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_347; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_348; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_349; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_350; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_351; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_352; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_353; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_354; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_355; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_356; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_357; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_358; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_359; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_360; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_361; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_362; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_363; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_364; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_365; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_366; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_367; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_368; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_369; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_370; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_371; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_372; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_373; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_374; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_375; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_376; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_377; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_378; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_379; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_380; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_381; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_382; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_383; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_384; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_385; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_386; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_387; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_388; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_389; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_390; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_391; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_392; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_393; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_394; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_395; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_396; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_397; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_398; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_399; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_400; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_401; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_402; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_403; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_404; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_405; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_406; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_407; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_408; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_409; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_410; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_411; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_412; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_413; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_414; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_415; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_416; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_417; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_418; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_419; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_420; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_421; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_422; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_423; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_424; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_425; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_426; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_427; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_428; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_429; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_430; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_431; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_432; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_433; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_434; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_435; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_436; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_437; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_438; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_439; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_440; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_441; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_442; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_443; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_444; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_445; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_446; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_447; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_448; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_449; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_450; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_451; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_452; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_453; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_454; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_455; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_456; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_457; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_458; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_459; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_460; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_461; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_462; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_463; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_464; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_465; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_466; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_467; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_468; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_469; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_470; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_471; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_472; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_473; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_474; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_475; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_476; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_477; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_478; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_479; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_480; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_481; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_482; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_483; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_484; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_485; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_486; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_487; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_488; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_489; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_490; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_491; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_492; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_493; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_494; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_495; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_496; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_497; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_498; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_499; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_500; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_501; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_502; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_503; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_504; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_505; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_506; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_507; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_508; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_509; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_510; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_511; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_512; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_513; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_514; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_515; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_516; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_517; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_518; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_519; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_520; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_521; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_522; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_523; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_524; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_525; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_526; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_527; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_528; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_529; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_530; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_531; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_532; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_533; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_534; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_535; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_536; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_537; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_538; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_539; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_540; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_541; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_542; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_543; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_544; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_545; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_546; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_547; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_548; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_549; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_550; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_551; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_552; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_553; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_554; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_555; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_556; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_557; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_558; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_559; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_560; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_561; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_562; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_563; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_564; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_565; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_566; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_567; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_568; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_569; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_570; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_571; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_572; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_573; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_574; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_575; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_576; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_577; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_578; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_579; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_580; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_581; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_582; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_583; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_584; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_585; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_586; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_587; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_588; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_589; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_590; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_591; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_592; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_593; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_594; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_595; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_596; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_597; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_598; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_599; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_600; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_601; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_602; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_603; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_604; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_605; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_606; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_607; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_608; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_609; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_610; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_611; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_612; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_613; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_614; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_615; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_616; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_617; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_618; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_619; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_620; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_621; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_622; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_623; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_624; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_625; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_626; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_627; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_628; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_629; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_630; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_631; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_632; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_633; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_634; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_635; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_636; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_637; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_638; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_639; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_640; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_641; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_642; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_643; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_644; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_645; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_646; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_647; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_648; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_649; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_650; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_651; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_652; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_653; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_654; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_655; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_656; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_657; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_658; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_659; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_660; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_661; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_662; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_663; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_664; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_665; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_666; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_667; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_668; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_669; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_670; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_671; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_672; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_673; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_674; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_675; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_676; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_677; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_678; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_679; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_680; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_681; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_682; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_683; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_684; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_685; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_686; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_687; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_688; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_689; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_690; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_691; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_692; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_693; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_694; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_695; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_696; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_697; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_698; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_699; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_700; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_701; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_702; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_703; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_704; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_705; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_706; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_707; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_708; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_709; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_710; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_711; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_712; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_713; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_714; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_715; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_716; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_717; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_718; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_719; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_720; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_721; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_722; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_723; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_724; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_725; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_726; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_727; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_728; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_729; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_730; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_731; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_732; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_733; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_734; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_735; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_736; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_737; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_738; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_739; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_740; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_741; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_742; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_743; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_744; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_745; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_746; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_747; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_748; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_749; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_750; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_751; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_752; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_753; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_754; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_755; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_756; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_757; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_758; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_759; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_760; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_761; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_762; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_763; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_764; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_765; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_766; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_767; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_768; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_769; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_770; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_771; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_772; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_773; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_774; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_775; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_776; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_777; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_778; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_779; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_780; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_781; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_782; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_783; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_784; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_785; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_786; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_787; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_788; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_789; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_790; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_791; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_792; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_793; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_794; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_795; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_796; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_797; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_798; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_799; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_800; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_801; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_802; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_803; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_804; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_805; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_806; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_807; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_808; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_809; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_810; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_811; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_812; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_813; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_814; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_815; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_816; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_817; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_818; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_819; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_820; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_821; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_822; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_823; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_824; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_825; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_826; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_827; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_828; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_829; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_830; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_831; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_832; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_833; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_834; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_835; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_836; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_837; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_838; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_839; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_840; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_841; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_842; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_843; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_844; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_845; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_846; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_847; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_848; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_849; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_850; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_851; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_852; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_853; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_854; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_855; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_856; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_857; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_858; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_859; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_860; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_861; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_862; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_863; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_864; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_865; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_866; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_867; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_868; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_869; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_870; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_871; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_872; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_873; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_874; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_875; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_876; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_877; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_878; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_879; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_880; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_881; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_882; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_883; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_884; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_885; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_886; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_887; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_888; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_889; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_890; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_891; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_892; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_893; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_894; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_895; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_896; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_897; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_898; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_899; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_900; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_901; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_902; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_903; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_904; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_905; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_906; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_907; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_908; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_909; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_910; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_911; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_912; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_913; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_914; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_915; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_916; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_917; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_918; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_919; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_920; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_921; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_922; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_923; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_924; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_925; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_926; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_927; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_928; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_929; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_930; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_931; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_932; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_933; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_934; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_935; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_936; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_937; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_938; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_939; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_940; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_941; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_942; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_943; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_944; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_945; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_946; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_947; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_948; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_949; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_950; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_951; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_952; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_953; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_954; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_955; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_956; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_957; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_958; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_959; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_960; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_961; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_962; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_963; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_964; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_965; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_966; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_967; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_968; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_969; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_970; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_971; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_972; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_973; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_974; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_975; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_976; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_977; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_978; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_979; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_980; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_981; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_982; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_983; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_984; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_985; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_986; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_987; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_988; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_989; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_990; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_991; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_992; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_993; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_994; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_995; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_996; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_997; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_998; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_999; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1000; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1001; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1002; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1003; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1004; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1005; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1006; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1007; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1008; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1009; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1010; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1011; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1012; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1013; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1014; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1015; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1016; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1017; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1018; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1019; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1020; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1021; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1022; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1023; // @[LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_0 = 10'h0 == io_wrAddr_0 ? 2'h0 : lvtReg_0; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1 = 10'h1 == io_wrAddr_0 ? 2'h0 : lvtReg_1; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2 = 10'h2 == io_wrAddr_0 ? 2'h0 : lvtReg_2; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_3 = 10'h3 == io_wrAddr_0 ? 2'h0 : lvtReg_3; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_4 = 10'h4 == io_wrAddr_0 ? 2'h0 : lvtReg_4; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_5 = 10'h5 == io_wrAddr_0 ? 2'h0 : lvtReg_5; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_6 = 10'h6 == io_wrAddr_0 ? 2'h0 : lvtReg_6; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_7 = 10'h7 == io_wrAddr_0 ? 2'h0 : lvtReg_7; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_8 = 10'h8 == io_wrAddr_0 ? 2'h0 : lvtReg_8; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_9 = 10'h9 == io_wrAddr_0 ? 2'h0 : lvtReg_9; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_10 = 10'ha == io_wrAddr_0 ? 2'h0 : lvtReg_10; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_11 = 10'hb == io_wrAddr_0 ? 2'h0 : lvtReg_11; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_12 = 10'hc == io_wrAddr_0 ? 2'h0 : lvtReg_12; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_13 = 10'hd == io_wrAddr_0 ? 2'h0 : lvtReg_13; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_14 = 10'he == io_wrAddr_0 ? 2'h0 : lvtReg_14; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_15 = 10'hf == io_wrAddr_0 ? 2'h0 : lvtReg_15; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_16 = 10'h10 == io_wrAddr_0 ? 2'h0 : lvtReg_16; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_17 = 10'h11 == io_wrAddr_0 ? 2'h0 : lvtReg_17; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_18 = 10'h12 == io_wrAddr_0 ? 2'h0 : lvtReg_18; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_19 = 10'h13 == io_wrAddr_0 ? 2'h0 : lvtReg_19; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_20 = 10'h14 == io_wrAddr_0 ? 2'h0 : lvtReg_20; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_21 = 10'h15 == io_wrAddr_0 ? 2'h0 : lvtReg_21; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_22 = 10'h16 == io_wrAddr_0 ? 2'h0 : lvtReg_22; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_23 = 10'h17 == io_wrAddr_0 ? 2'h0 : lvtReg_23; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_24 = 10'h18 == io_wrAddr_0 ? 2'h0 : lvtReg_24; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_25 = 10'h19 == io_wrAddr_0 ? 2'h0 : lvtReg_25; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_26 = 10'h1a == io_wrAddr_0 ? 2'h0 : lvtReg_26; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_27 = 10'h1b == io_wrAddr_0 ? 2'h0 : lvtReg_27; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_28 = 10'h1c == io_wrAddr_0 ? 2'h0 : lvtReg_28; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_29 = 10'h1d == io_wrAddr_0 ? 2'h0 : lvtReg_29; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_30 = 10'h1e == io_wrAddr_0 ? 2'h0 : lvtReg_30; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_31 = 10'h1f == io_wrAddr_0 ? 2'h0 : lvtReg_31; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_32 = 10'h20 == io_wrAddr_0 ? 2'h0 : lvtReg_32; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_33 = 10'h21 == io_wrAddr_0 ? 2'h0 : lvtReg_33; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_34 = 10'h22 == io_wrAddr_0 ? 2'h0 : lvtReg_34; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_35 = 10'h23 == io_wrAddr_0 ? 2'h0 : lvtReg_35; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_36 = 10'h24 == io_wrAddr_0 ? 2'h0 : lvtReg_36; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_37 = 10'h25 == io_wrAddr_0 ? 2'h0 : lvtReg_37; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_38 = 10'h26 == io_wrAddr_0 ? 2'h0 : lvtReg_38; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_39 = 10'h27 == io_wrAddr_0 ? 2'h0 : lvtReg_39; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_40 = 10'h28 == io_wrAddr_0 ? 2'h0 : lvtReg_40; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_41 = 10'h29 == io_wrAddr_0 ? 2'h0 : lvtReg_41; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_42 = 10'h2a == io_wrAddr_0 ? 2'h0 : lvtReg_42; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_43 = 10'h2b == io_wrAddr_0 ? 2'h0 : lvtReg_43; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_44 = 10'h2c == io_wrAddr_0 ? 2'h0 : lvtReg_44; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_45 = 10'h2d == io_wrAddr_0 ? 2'h0 : lvtReg_45; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_46 = 10'h2e == io_wrAddr_0 ? 2'h0 : lvtReg_46; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_47 = 10'h2f == io_wrAddr_0 ? 2'h0 : lvtReg_47; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_48 = 10'h30 == io_wrAddr_0 ? 2'h0 : lvtReg_48; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_49 = 10'h31 == io_wrAddr_0 ? 2'h0 : lvtReg_49; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_50 = 10'h32 == io_wrAddr_0 ? 2'h0 : lvtReg_50; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_51 = 10'h33 == io_wrAddr_0 ? 2'h0 : lvtReg_51; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_52 = 10'h34 == io_wrAddr_0 ? 2'h0 : lvtReg_52; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_53 = 10'h35 == io_wrAddr_0 ? 2'h0 : lvtReg_53; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_54 = 10'h36 == io_wrAddr_0 ? 2'h0 : lvtReg_54; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_55 = 10'h37 == io_wrAddr_0 ? 2'h0 : lvtReg_55; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_56 = 10'h38 == io_wrAddr_0 ? 2'h0 : lvtReg_56; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_57 = 10'h39 == io_wrAddr_0 ? 2'h0 : lvtReg_57; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_58 = 10'h3a == io_wrAddr_0 ? 2'h0 : lvtReg_58; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_59 = 10'h3b == io_wrAddr_0 ? 2'h0 : lvtReg_59; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_60 = 10'h3c == io_wrAddr_0 ? 2'h0 : lvtReg_60; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_61 = 10'h3d == io_wrAddr_0 ? 2'h0 : lvtReg_61; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_62 = 10'h3e == io_wrAddr_0 ? 2'h0 : lvtReg_62; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_63 = 10'h3f == io_wrAddr_0 ? 2'h0 : lvtReg_63; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_64 = 10'h40 == io_wrAddr_0 ? 2'h0 : lvtReg_64; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_65 = 10'h41 == io_wrAddr_0 ? 2'h0 : lvtReg_65; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_66 = 10'h42 == io_wrAddr_0 ? 2'h0 : lvtReg_66; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_67 = 10'h43 == io_wrAddr_0 ? 2'h0 : lvtReg_67; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_68 = 10'h44 == io_wrAddr_0 ? 2'h0 : lvtReg_68; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_69 = 10'h45 == io_wrAddr_0 ? 2'h0 : lvtReg_69; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_70 = 10'h46 == io_wrAddr_0 ? 2'h0 : lvtReg_70; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_71 = 10'h47 == io_wrAddr_0 ? 2'h0 : lvtReg_71; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_72 = 10'h48 == io_wrAddr_0 ? 2'h0 : lvtReg_72; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_73 = 10'h49 == io_wrAddr_0 ? 2'h0 : lvtReg_73; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_74 = 10'h4a == io_wrAddr_0 ? 2'h0 : lvtReg_74; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_75 = 10'h4b == io_wrAddr_0 ? 2'h0 : lvtReg_75; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_76 = 10'h4c == io_wrAddr_0 ? 2'h0 : lvtReg_76; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_77 = 10'h4d == io_wrAddr_0 ? 2'h0 : lvtReg_77; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_78 = 10'h4e == io_wrAddr_0 ? 2'h0 : lvtReg_78; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_79 = 10'h4f == io_wrAddr_0 ? 2'h0 : lvtReg_79; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_80 = 10'h50 == io_wrAddr_0 ? 2'h0 : lvtReg_80; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_81 = 10'h51 == io_wrAddr_0 ? 2'h0 : lvtReg_81; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_82 = 10'h52 == io_wrAddr_0 ? 2'h0 : lvtReg_82; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_83 = 10'h53 == io_wrAddr_0 ? 2'h0 : lvtReg_83; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_84 = 10'h54 == io_wrAddr_0 ? 2'h0 : lvtReg_84; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_85 = 10'h55 == io_wrAddr_0 ? 2'h0 : lvtReg_85; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_86 = 10'h56 == io_wrAddr_0 ? 2'h0 : lvtReg_86; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_87 = 10'h57 == io_wrAddr_0 ? 2'h0 : lvtReg_87; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_88 = 10'h58 == io_wrAddr_0 ? 2'h0 : lvtReg_88; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_89 = 10'h59 == io_wrAddr_0 ? 2'h0 : lvtReg_89; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_90 = 10'h5a == io_wrAddr_0 ? 2'h0 : lvtReg_90; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_91 = 10'h5b == io_wrAddr_0 ? 2'h0 : lvtReg_91; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_92 = 10'h5c == io_wrAddr_0 ? 2'h0 : lvtReg_92; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_93 = 10'h5d == io_wrAddr_0 ? 2'h0 : lvtReg_93; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_94 = 10'h5e == io_wrAddr_0 ? 2'h0 : lvtReg_94; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_95 = 10'h5f == io_wrAddr_0 ? 2'h0 : lvtReg_95; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_96 = 10'h60 == io_wrAddr_0 ? 2'h0 : lvtReg_96; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_97 = 10'h61 == io_wrAddr_0 ? 2'h0 : lvtReg_97; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_98 = 10'h62 == io_wrAddr_0 ? 2'h0 : lvtReg_98; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_99 = 10'h63 == io_wrAddr_0 ? 2'h0 : lvtReg_99; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_100 = 10'h64 == io_wrAddr_0 ? 2'h0 : lvtReg_100; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_101 = 10'h65 == io_wrAddr_0 ? 2'h0 : lvtReg_101; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_102 = 10'h66 == io_wrAddr_0 ? 2'h0 : lvtReg_102; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_103 = 10'h67 == io_wrAddr_0 ? 2'h0 : lvtReg_103; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_104 = 10'h68 == io_wrAddr_0 ? 2'h0 : lvtReg_104; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_105 = 10'h69 == io_wrAddr_0 ? 2'h0 : lvtReg_105; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_106 = 10'h6a == io_wrAddr_0 ? 2'h0 : lvtReg_106; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_107 = 10'h6b == io_wrAddr_0 ? 2'h0 : lvtReg_107; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_108 = 10'h6c == io_wrAddr_0 ? 2'h0 : lvtReg_108; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_109 = 10'h6d == io_wrAddr_0 ? 2'h0 : lvtReg_109; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_110 = 10'h6e == io_wrAddr_0 ? 2'h0 : lvtReg_110; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_111 = 10'h6f == io_wrAddr_0 ? 2'h0 : lvtReg_111; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_112 = 10'h70 == io_wrAddr_0 ? 2'h0 : lvtReg_112; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_113 = 10'h71 == io_wrAddr_0 ? 2'h0 : lvtReg_113; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_114 = 10'h72 == io_wrAddr_0 ? 2'h0 : lvtReg_114; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_115 = 10'h73 == io_wrAddr_0 ? 2'h0 : lvtReg_115; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_116 = 10'h74 == io_wrAddr_0 ? 2'h0 : lvtReg_116; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_117 = 10'h75 == io_wrAddr_0 ? 2'h0 : lvtReg_117; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_118 = 10'h76 == io_wrAddr_0 ? 2'h0 : lvtReg_118; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_119 = 10'h77 == io_wrAddr_0 ? 2'h0 : lvtReg_119; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_120 = 10'h78 == io_wrAddr_0 ? 2'h0 : lvtReg_120; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_121 = 10'h79 == io_wrAddr_0 ? 2'h0 : lvtReg_121; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_122 = 10'h7a == io_wrAddr_0 ? 2'h0 : lvtReg_122; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_123 = 10'h7b == io_wrAddr_0 ? 2'h0 : lvtReg_123; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_124 = 10'h7c == io_wrAddr_0 ? 2'h0 : lvtReg_124; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_125 = 10'h7d == io_wrAddr_0 ? 2'h0 : lvtReg_125; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_126 = 10'h7e == io_wrAddr_0 ? 2'h0 : lvtReg_126; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_127 = 10'h7f == io_wrAddr_0 ? 2'h0 : lvtReg_127; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_128 = 10'h80 == io_wrAddr_0 ? 2'h0 : lvtReg_128; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_129 = 10'h81 == io_wrAddr_0 ? 2'h0 : lvtReg_129; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_130 = 10'h82 == io_wrAddr_0 ? 2'h0 : lvtReg_130; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_131 = 10'h83 == io_wrAddr_0 ? 2'h0 : lvtReg_131; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_132 = 10'h84 == io_wrAddr_0 ? 2'h0 : lvtReg_132; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_133 = 10'h85 == io_wrAddr_0 ? 2'h0 : lvtReg_133; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_134 = 10'h86 == io_wrAddr_0 ? 2'h0 : lvtReg_134; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_135 = 10'h87 == io_wrAddr_0 ? 2'h0 : lvtReg_135; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_136 = 10'h88 == io_wrAddr_0 ? 2'h0 : lvtReg_136; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_137 = 10'h89 == io_wrAddr_0 ? 2'h0 : lvtReg_137; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_138 = 10'h8a == io_wrAddr_0 ? 2'h0 : lvtReg_138; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_139 = 10'h8b == io_wrAddr_0 ? 2'h0 : lvtReg_139; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_140 = 10'h8c == io_wrAddr_0 ? 2'h0 : lvtReg_140; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_141 = 10'h8d == io_wrAddr_0 ? 2'h0 : lvtReg_141; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_142 = 10'h8e == io_wrAddr_0 ? 2'h0 : lvtReg_142; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_143 = 10'h8f == io_wrAddr_0 ? 2'h0 : lvtReg_143; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_144 = 10'h90 == io_wrAddr_0 ? 2'h0 : lvtReg_144; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_145 = 10'h91 == io_wrAddr_0 ? 2'h0 : lvtReg_145; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_146 = 10'h92 == io_wrAddr_0 ? 2'h0 : lvtReg_146; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_147 = 10'h93 == io_wrAddr_0 ? 2'h0 : lvtReg_147; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_148 = 10'h94 == io_wrAddr_0 ? 2'h0 : lvtReg_148; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_149 = 10'h95 == io_wrAddr_0 ? 2'h0 : lvtReg_149; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_150 = 10'h96 == io_wrAddr_0 ? 2'h0 : lvtReg_150; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_151 = 10'h97 == io_wrAddr_0 ? 2'h0 : lvtReg_151; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_152 = 10'h98 == io_wrAddr_0 ? 2'h0 : lvtReg_152; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_153 = 10'h99 == io_wrAddr_0 ? 2'h0 : lvtReg_153; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_154 = 10'h9a == io_wrAddr_0 ? 2'h0 : lvtReg_154; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_155 = 10'h9b == io_wrAddr_0 ? 2'h0 : lvtReg_155; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_156 = 10'h9c == io_wrAddr_0 ? 2'h0 : lvtReg_156; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_157 = 10'h9d == io_wrAddr_0 ? 2'h0 : lvtReg_157; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_158 = 10'h9e == io_wrAddr_0 ? 2'h0 : lvtReg_158; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_159 = 10'h9f == io_wrAddr_0 ? 2'h0 : lvtReg_159; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_160 = 10'ha0 == io_wrAddr_0 ? 2'h0 : lvtReg_160; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_161 = 10'ha1 == io_wrAddr_0 ? 2'h0 : lvtReg_161; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_162 = 10'ha2 == io_wrAddr_0 ? 2'h0 : lvtReg_162; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_163 = 10'ha3 == io_wrAddr_0 ? 2'h0 : lvtReg_163; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_164 = 10'ha4 == io_wrAddr_0 ? 2'h0 : lvtReg_164; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_165 = 10'ha5 == io_wrAddr_0 ? 2'h0 : lvtReg_165; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_166 = 10'ha6 == io_wrAddr_0 ? 2'h0 : lvtReg_166; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_167 = 10'ha7 == io_wrAddr_0 ? 2'h0 : lvtReg_167; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_168 = 10'ha8 == io_wrAddr_0 ? 2'h0 : lvtReg_168; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_169 = 10'ha9 == io_wrAddr_0 ? 2'h0 : lvtReg_169; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_170 = 10'haa == io_wrAddr_0 ? 2'h0 : lvtReg_170; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_171 = 10'hab == io_wrAddr_0 ? 2'h0 : lvtReg_171; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_172 = 10'hac == io_wrAddr_0 ? 2'h0 : lvtReg_172; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_173 = 10'had == io_wrAddr_0 ? 2'h0 : lvtReg_173; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_174 = 10'hae == io_wrAddr_0 ? 2'h0 : lvtReg_174; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_175 = 10'haf == io_wrAddr_0 ? 2'h0 : lvtReg_175; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_176 = 10'hb0 == io_wrAddr_0 ? 2'h0 : lvtReg_176; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_177 = 10'hb1 == io_wrAddr_0 ? 2'h0 : lvtReg_177; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_178 = 10'hb2 == io_wrAddr_0 ? 2'h0 : lvtReg_178; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_179 = 10'hb3 == io_wrAddr_0 ? 2'h0 : lvtReg_179; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_180 = 10'hb4 == io_wrAddr_0 ? 2'h0 : lvtReg_180; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_181 = 10'hb5 == io_wrAddr_0 ? 2'h0 : lvtReg_181; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_182 = 10'hb6 == io_wrAddr_0 ? 2'h0 : lvtReg_182; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_183 = 10'hb7 == io_wrAddr_0 ? 2'h0 : lvtReg_183; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_184 = 10'hb8 == io_wrAddr_0 ? 2'h0 : lvtReg_184; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_185 = 10'hb9 == io_wrAddr_0 ? 2'h0 : lvtReg_185; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_186 = 10'hba == io_wrAddr_0 ? 2'h0 : lvtReg_186; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_187 = 10'hbb == io_wrAddr_0 ? 2'h0 : lvtReg_187; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_188 = 10'hbc == io_wrAddr_0 ? 2'h0 : lvtReg_188; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_189 = 10'hbd == io_wrAddr_0 ? 2'h0 : lvtReg_189; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_190 = 10'hbe == io_wrAddr_0 ? 2'h0 : lvtReg_190; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_191 = 10'hbf == io_wrAddr_0 ? 2'h0 : lvtReg_191; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_192 = 10'hc0 == io_wrAddr_0 ? 2'h0 : lvtReg_192; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_193 = 10'hc1 == io_wrAddr_0 ? 2'h0 : lvtReg_193; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_194 = 10'hc2 == io_wrAddr_0 ? 2'h0 : lvtReg_194; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_195 = 10'hc3 == io_wrAddr_0 ? 2'h0 : lvtReg_195; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_196 = 10'hc4 == io_wrAddr_0 ? 2'h0 : lvtReg_196; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_197 = 10'hc5 == io_wrAddr_0 ? 2'h0 : lvtReg_197; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_198 = 10'hc6 == io_wrAddr_0 ? 2'h0 : lvtReg_198; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_199 = 10'hc7 == io_wrAddr_0 ? 2'h0 : lvtReg_199; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_200 = 10'hc8 == io_wrAddr_0 ? 2'h0 : lvtReg_200; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_201 = 10'hc9 == io_wrAddr_0 ? 2'h0 : lvtReg_201; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_202 = 10'hca == io_wrAddr_0 ? 2'h0 : lvtReg_202; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_203 = 10'hcb == io_wrAddr_0 ? 2'h0 : lvtReg_203; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_204 = 10'hcc == io_wrAddr_0 ? 2'h0 : lvtReg_204; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_205 = 10'hcd == io_wrAddr_0 ? 2'h0 : lvtReg_205; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_206 = 10'hce == io_wrAddr_0 ? 2'h0 : lvtReg_206; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_207 = 10'hcf == io_wrAddr_0 ? 2'h0 : lvtReg_207; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_208 = 10'hd0 == io_wrAddr_0 ? 2'h0 : lvtReg_208; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_209 = 10'hd1 == io_wrAddr_0 ? 2'h0 : lvtReg_209; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_210 = 10'hd2 == io_wrAddr_0 ? 2'h0 : lvtReg_210; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_211 = 10'hd3 == io_wrAddr_0 ? 2'h0 : lvtReg_211; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_212 = 10'hd4 == io_wrAddr_0 ? 2'h0 : lvtReg_212; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_213 = 10'hd5 == io_wrAddr_0 ? 2'h0 : lvtReg_213; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_214 = 10'hd6 == io_wrAddr_0 ? 2'h0 : lvtReg_214; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_215 = 10'hd7 == io_wrAddr_0 ? 2'h0 : lvtReg_215; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_216 = 10'hd8 == io_wrAddr_0 ? 2'h0 : lvtReg_216; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_217 = 10'hd9 == io_wrAddr_0 ? 2'h0 : lvtReg_217; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_218 = 10'hda == io_wrAddr_0 ? 2'h0 : lvtReg_218; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_219 = 10'hdb == io_wrAddr_0 ? 2'h0 : lvtReg_219; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_220 = 10'hdc == io_wrAddr_0 ? 2'h0 : lvtReg_220; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_221 = 10'hdd == io_wrAddr_0 ? 2'h0 : lvtReg_221; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_222 = 10'hde == io_wrAddr_0 ? 2'h0 : lvtReg_222; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_223 = 10'hdf == io_wrAddr_0 ? 2'h0 : lvtReg_223; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_224 = 10'he0 == io_wrAddr_0 ? 2'h0 : lvtReg_224; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_225 = 10'he1 == io_wrAddr_0 ? 2'h0 : lvtReg_225; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_226 = 10'he2 == io_wrAddr_0 ? 2'h0 : lvtReg_226; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_227 = 10'he3 == io_wrAddr_0 ? 2'h0 : lvtReg_227; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_228 = 10'he4 == io_wrAddr_0 ? 2'h0 : lvtReg_228; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_229 = 10'he5 == io_wrAddr_0 ? 2'h0 : lvtReg_229; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_230 = 10'he6 == io_wrAddr_0 ? 2'h0 : lvtReg_230; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_231 = 10'he7 == io_wrAddr_0 ? 2'h0 : lvtReg_231; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_232 = 10'he8 == io_wrAddr_0 ? 2'h0 : lvtReg_232; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_233 = 10'he9 == io_wrAddr_0 ? 2'h0 : lvtReg_233; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_234 = 10'hea == io_wrAddr_0 ? 2'h0 : lvtReg_234; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_235 = 10'heb == io_wrAddr_0 ? 2'h0 : lvtReg_235; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_236 = 10'hec == io_wrAddr_0 ? 2'h0 : lvtReg_236; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_237 = 10'hed == io_wrAddr_0 ? 2'h0 : lvtReg_237; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_238 = 10'hee == io_wrAddr_0 ? 2'h0 : lvtReg_238; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_239 = 10'hef == io_wrAddr_0 ? 2'h0 : lvtReg_239; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_240 = 10'hf0 == io_wrAddr_0 ? 2'h0 : lvtReg_240; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_241 = 10'hf1 == io_wrAddr_0 ? 2'h0 : lvtReg_241; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_242 = 10'hf2 == io_wrAddr_0 ? 2'h0 : lvtReg_242; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_243 = 10'hf3 == io_wrAddr_0 ? 2'h0 : lvtReg_243; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_244 = 10'hf4 == io_wrAddr_0 ? 2'h0 : lvtReg_244; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_245 = 10'hf5 == io_wrAddr_0 ? 2'h0 : lvtReg_245; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_246 = 10'hf6 == io_wrAddr_0 ? 2'h0 : lvtReg_246; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_247 = 10'hf7 == io_wrAddr_0 ? 2'h0 : lvtReg_247; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_248 = 10'hf8 == io_wrAddr_0 ? 2'h0 : lvtReg_248; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_249 = 10'hf9 == io_wrAddr_0 ? 2'h0 : lvtReg_249; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_250 = 10'hfa == io_wrAddr_0 ? 2'h0 : lvtReg_250; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_251 = 10'hfb == io_wrAddr_0 ? 2'h0 : lvtReg_251; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_252 = 10'hfc == io_wrAddr_0 ? 2'h0 : lvtReg_252; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_253 = 10'hfd == io_wrAddr_0 ? 2'h0 : lvtReg_253; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_254 = 10'hfe == io_wrAddr_0 ? 2'h0 : lvtReg_254; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_255 = 10'hff == io_wrAddr_0 ? 2'h0 : lvtReg_255; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_256 = 10'h100 == io_wrAddr_0 ? 2'h0 : lvtReg_256; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_257 = 10'h101 == io_wrAddr_0 ? 2'h0 : lvtReg_257; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_258 = 10'h102 == io_wrAddr_0 ? 2'h0 : lvtReg_258; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_259 = 10'h103 == io_wrAddr_0 ? 2'h0 : lvtReg_259; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_260 = 10'h104 == io_wrAddr_0 ? 2'h0 : lvtReg_260; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_261 = 10'h105 == io_wrAddr_0 ? 2'h0 : lvtReg_261; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_262 = 10'h106 == io_wrAddr_0 ? 2'h0 : lvtReg_262; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_263 = 10'h107 == io_wrAddr_0 ? 2'h0 : lvtReg_263; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_264 = 10'h108 == io_wrAddr_0 ? 2'h0 : lvtReg_264; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_265 = 10'h109 == io_wrAddr_0 ? 2'h0 : lvtReg_265; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_266 = 10'h10a == io_wrAddr_0 ? 2'h0 : lvtReg_266; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_267 = 10'h10b == io_wrAddr_0 ? 2'h0 : lvtReg_267; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_268 = 10'h10c == io_wrAddr_0 ? 2'h0 : lvtReg_268; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_269 = 10'h10d == io_wrAddr_0 ? 2'h0 : lvtReg_269; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_270 = 10'h10e == io_wrAddr_0 ? 2'h0 : lvtReg_270; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_271 = 10'h10f == io_wrAddr_0 ? 2'h0 : lvtReg_271; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_272 = 10'h110 == io_wrAddr_0 ? 2'h0 : lvtReg_272; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_273 = 10'h111 == io_wrAddr_0 ? 2'h0 : lvtReg_273; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_274 = 10'h112 == io_wrAddr_0 ? 2'h0 : lvtReg_274; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_275 = 10'h113 == io_wrAddr_0 ? 2'h0 : lvtReg_275; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_276 = 10'h114 == io_wrAddr_0 ? 2'h0 : lvtReg_276; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_277 = 10'h115 == io_wrAddr_0 ? 2'h0 : lvtReg_277; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_278 = 10'h116 == io_wrAddr_0 ? 2'h0 : lvtReg_278; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_279 = 10'h117 == io_wrAddr_0 ? 2'h0 : lvtReg_279; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_280 = 10'h118 == io_wrAddr_0 ? 2'h0 : lvtReg_280; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_281 = 10'h119 == io_wrAddr_0 ? 2'h0 : lvtReg_281; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_282 = 10'h11a == io_wrAddr_0 ? 2'h0 : lvtReg_282; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_283 = 10'h11b == io_wrAddr_0 ? 2'h0 : lvtReg_283; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_284 = 10'h11c == io_wrAddr_0 ? 2'h0 : lvtReg_284; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_285 = 10'h11d == io_wrAddr_0 ? 2'h0 : lvtReg_285; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_286 = 10'h11e == io_wrAddr_0 ? 2'h0 : lvtReg_286; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_287 = 10'h11f == io_wrAddr_0 ? 2'h0 : lvtReg_287; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_288 = 10'h120 == io_wrAddr_0 ? 2'h0 : lvtReg_288; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_289 = 10'h121 == io_wrAddr_0 ? 2'h0 : lvtReg_289; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_290 = 10'h122 == io_wrAddr_0 ? 2'h0 : lvtReg_290; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_291 = 10'h123 == io_wrAddr_0 ? 2'h0 : lvtReg_291; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_292 = 10'h124 == io_wrAddr_0 ? 2'h0 : lvtReg_292; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_293 = 10'h125 == io_wrAddr_0 ? 2'h0 : lvtReg_293; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_294 = 10'h126 == io_wrAddr_0 ? 2'h0 : lvtReg_294; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_295 = 10'h127 == io_wrAddr_0 ? 2'h0 : lvtReg_295; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_296 = 10'h128 == io_wrAddr_0 ? 2'h0 : lvtReg_296; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_297 = 10'h129 == io_wrAddr_0 ? 2'h0 : lvtReg_297; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_298 = 10'h12a == io_wrAddr_0 ? 2'h0 : lvtReg_298; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_299 = 10'h12b == io_wrAddr_0 ? 2'h0 : lvtReg_299; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_300 = 10'h12c == io_wrAddr_0 ? 2'h0 : lvtReg_300; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_301 = 10'h12d == io_wrAddr_0 ? 2'h0 : lvtReg_301; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_302 = 10'h12e == io_wrAddr_0 ? 2'h0 : lvtReg_302; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_303 = 10'h12f == io_wrAddr_0 ? 2'h0 : lvtReg_303; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_304 = 10'h130 == io_wrAddr_0 ? 2'h0 : lvtReg_304; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_305 = 10'h131 == io_wrAddr_0 ? 2'h0 : lvtReg_305; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_306 = 10'h132 == io_wrAddr_0 ? 2'h0 : lvtReg_306; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_307 = 10'h133 == io_wrAddr_0 ? 2'h0 : lvtReg_307; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_308 = 10'h134 == io_wrAddr_0 ? 2'h0 : lvtReg_308; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_309 = 10'h135 == io_wrAddr_0 ? 2'h0 : lvtReg_309; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_310 = 10'h136 == io_wrAddr_0 ? 2'h0 : lvtReg_310; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_311 = 10'h137 == io_wrAddr_0 ? 2'h0 : lvtReg_311; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_312 = 10'h138 == io_wrAddr_0 ? 2'h0 : lvtReg_312; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_313 = 10'h139 == io_wrAddr_0 ? 2'h0 : lvtReg_313; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_314 = 10'h13a == io_wrAddr_0 ? 2'h0 : lvtReg_314; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_315 = 10'h13b == io_wrAddr_0 ? 2'h0 : lvtReg_315; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_316 = 10'h13c == io_wrAddr_0 ? 2'h0 : lvtReg_316; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_317 = 10'h13d == io_wrAddr_0 ? 2'h0 : lvtReg_317; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_318 = 10'h13e == io_wrAddr_0 ? 2'h0 : lvtReg_318; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_319 = 10'h13f == io_wrAddr_0 ? 2'h0 : lvtReg_319; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_320 = 10'h140 == io_wrAddr_0 ? 2'h0 : lvtReg_320; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_321 = 10'h141 == io_wrAddr_0 ? 2'h0 : lvtReg_321; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_322 = 10'h142 == io_wrAddr_0 ? 2'h0 : lvtReg_322; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_323 = 10'h143 == io_wrAddr_0 ? 2'h0 : lvtReg_323; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_324 = 10'h144 == io_wrAddr_0 ? 2'h0 : lvtReg_324; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_325 = 10'h145 == io_wrAddr_0 ? 2'h0 : lvtReg_325; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_326 = 10'h146 == io_wrAddr_0 ? 2'h0 : lvtReg_326; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_327 = 10'h147 == io_wrAddr_0 ? 2'h0 : lvtReg_327; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_328 = 10'h148 == io_wrAddr_0 ? 2'h0 : lvtReg_328; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_329 = 10'h149 == io_wrAddr_0 ? 2'h0 : lvtReg_329; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_330 = 10'h14a == io_wrAddr_0 ? 2'h0 : lvtReg_330; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_331 = 10'h14b == io_wrAddr_0 ? 2'h0 : lvtReg_331; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_332 = 10'h14c == io_wrAddr_0 ? 2'h0 : lvtReg_332; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_333 = 10'h14d == io_wrAddr_0 ? 2'h0 : lvtReg_333; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_334 = 10'h14e == io_wrAddr_0 ? 2'h0 : lvtReg_334; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_335 = 10'h14f == io_wrAddr_0 ? 2'h0 : lvtReg_335; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_336 = 10'h150 == io_wrAddr_0 ? 2'h0 : lvtReg_336; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_337 = 10'h151 == io_wrAddr_0 ? 2'h0 : lvtReg_337; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_338 = 10'h152 == io_wrAddr_0 ? 2'h0 : lvtReg_338; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_339 = 10'h153 == io_wrAddr_0 ? 2'h0 : lvtReg_339; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_340 = 10'h154 == io_wrAddr_0 ? 2'h0 : lvtReg_340; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_341 = 10'h155 == io_wrAddr_0 ? 2'h0 : lvtReg_341; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_342 = 10'h156 == io_wrAddr_0 ? 2'h0 : lvtReg_342; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_343 = 10'h157 == io_wrAddr_0 ? 2'h0 : lvtReg_343; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_344 = 10'h158 == io_wrAddr_0 ? 2'h0 : lvtReg_344; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_345 = 10'h159 == io_wrAddr_0 ? 2'h0 : lvtReg_345; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_346 = 10'h15a == io_wrAddr_0 ? 2'h0 : lvtReg_346; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_347 = 10'h15b == io_wrAddr_0 ? 2'h0 : lvtReg_347; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_348 = 10'h15c == io_wrAddr_0 ? 2'h0 : lvtReg_348; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_349 = 10'h15d == io_wrAddr_0 ? 2'h0 : lvtReg_349; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_350 = 10'h15e == io_wrAddr_0 ? 2'h0 : lvtReg_350; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_351 = 10'h15f == io_wrAddr_0 ? 2'h0 : lvtReg_351; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_352 = 10'h160 == io_wrAddr_0 ? 2'h0 : lvtReg_352; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_353 = 10'h161 == io_wrAddr_0 ? 2'h0 : lvtReg_353; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_354 = 10'h162 == io_wrAddr_0 ? 2'h0 : lvtReg_354; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_355 = 10'h163 == io_wrAddr_0 ? 2'h0 : lvtReg_355; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_356 = 10'h164 == io_wrAddr_0 ? 2'h0 : lvtReg_356; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_357 = 10'h165 == io_wrAddr_0 ? 2'h0 : lvtReg_357; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_358 = 10'h166 == io_wrAddr_0 ? 2'h0 : lvtReg_358; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_359 = 10'h167 == io_wrAddr_0 ? 2'h0 : lvtReg_359; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_360 = 10'h168 == io_wrAddr_0 ? 2'h0 : lvtReg_360; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_361 = 10'h169 == io_wrAddr_0 ? 2'h0 : lvtReg_361; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_362 = 10'h16a == io_wrAddr_0 ? 2'h0 : lvtReg_362; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_363 = 10'h16b == io_wrAddr_0 ? 2'h0 : lvtReg_363; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_364 = 10'h16c == io_wrAddr_0 ? 2'h0 : lvtReg_364; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_365 = 10'h16d == io_wrAddr_0 ? 2'h0 : lvtReg_365; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_366 = 10'h16e == io_wrAddr_0 ? 2'h0 : lvtReg_366; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_367 = 10'h16f == io_wrAddr_0 ? 2'h0 : lvtReg_367; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_368 = 10'h170 == io_wrAddr_0 ? 2'h0 : lvtReg_368; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_369 = 10'h171 == io_wrAddr_0 ? 2'h0 : lvtReg_369; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_370 = 10'h172 == io_wrAddr_0 ? 2'h0 : lvtReg_370; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_371 = 10'h173 == io_wrAddr_0 ? 2'h0 : lvtReg_371; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_372 = 10'h174 == io_wrAddr_0 ? 2'h0 : lvtReg_372; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_373 = 10'h175 == io_wrAddr_0 ? 2'h0 : lvtReg_373; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_374 = 10'h176 == io_wrAddr_0 ? 2'h0 : lvtReg_374; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_375 = 10'h177 == io_wrAddr_0 ? 2'h0 : lvtReg_375; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_376 = 10'h178 == io_wrAddr_0 ? 2'h0 : lvtReg_376; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_377 = 10'h179 == io_wrAddr_0 ? 2'h0 : lvtReg_377; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_378 = 10'h17a == io_wrAddr_0 ? 2'h0 : lvtReg_378; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_379 = 10'h17b == io_wrAddr_0 ? 2'h0 : lvtReg_379; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_380 = 10'h17c == io_wrAddr_0 ? 2'h0 : lvtReg_380; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_381 = 10'h17d == io_wrAddr_0 ? 2'h0 : lvtReg_381; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_382 = 10'h17e == io_wrAddr_0 ? 2'h0 : lvtReg_382; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_383 = 10'h17f == io_wrAddr_0 ? 2'h0 : lvtReg_383; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_384 = 10'h180 == io_wrAddr_0 ? 2'h0 : lvtReg_384; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_385 = 10'h181 == io_wrAddr_0 ? 2'h0 : lvtReg_385; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_386 = 10'h182 == io_wrAddr_0 ? 2'h0 : lvtReg_386; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_387 = 10'h183 == io_wrAddr_0 ? 2'h0 : lvtReg_387; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_388 = 10'h184 == io_wrAddr_0 ? 2'h0 : lvtReg_388; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_389 = 10'h185 == io_wrAddr_0 ? 2'h0 : lvtReg_389; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_390 = 10'h186 == io_wrAddr_0 ? 2'h0 : lvtReg_390; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_391 = 10'h187 == io_wrAddr_0 ? 2'h0 : lvtReg_391; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_392 = 10'h188 == io_wrAddr_0 ? 2'h0 : lvtReg_392; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_393 = 10'h189 == io_wrAddr_0 ? 2'h0 : lvtReg_393; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_394 = 10'h18a == io_wrAddr_0 ? 2'h0 : lvtReg_394; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_395 = 10'h18b == io_wrAddr_0 ? 2'h0 : lvtReg_395; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_396 = 10'h18c == io_wrAddr_0 ? 2'h0 : lvtReg_396; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_397 = 10'h18d == io_wrAddr_0 ? 2'h0 : lvtReg_397; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_398 = 10'h18e == io_wrAddr_0 ? 2'h0 : lvtReg_398; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_399 = 10'h18f == io_wrAddr_0 ? 2'h0 : lvtReg_399; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_400 = 10'h190 == io_wrAddr_0 ? 2'h0 : lvtReg_400; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_401 = 10'h191 == io_wrAddr_0 ? 2'h0 : lvtReg_401; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_402 = 10'h192 == io_wrAddr_0 ? 2'h0 : lvtReg_402; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_403 = 10'h193 == io_wrAddr_0 ? 2'h0 : lvtReg_403; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_404 = 10'h194 == io_wrAddr_0 ? 2'h0 : lvtReg_404; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_405 = 10'h195 == io_wrAddr_0 ? 2'h0 : lvtReg_405; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_406 = 10'h196 == io_wrAddr_0 ? 2'h0 : lvtReg_406; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_407 = 10'h197 == io_wrAddr_0 ? 2'h0 : lvtReg_407; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_408 = 10'h198 == io_wrAddr_0 ? 2'h0 : lvtReg_408; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_409 = 10'h199 == io_wrAddr_0 ? 2'h0 : lvtReg_409; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_410 = 10'h19a == io_wrAddr_0 ? 2'h0 : lvtReg_410; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_411 = 10'h19b == io_wrAddr_0 ? 2'h0 : lvtReg_411; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_412 = 10'h19c == io_wrAddr_0 ? 2'h0 : lvtReg_412; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_413 = 10'h19d == io_wrAddr_0 ? 2'h0 : lvtReg_413; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_414 = 10'h19e == io_wrAddr_0 ? 2'h0 : lvtReg_414; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_415 = 10'h19f == io_wrAddr_0 ? 2'h0 : lvtReg_415; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_416 = 10'h1a0 == io_wrAddr_0 ? 2'h0 : lvtReg_416; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_417 = 10'h1a1 == io_wrAddr_0 ? 2'h0 : lvtReg_417; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_418 = 10'h1a2 == io_wrAddr_0 ? 2'h0 : lvtReg_418; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_419 = 10'h1a3 == io_wrAddr_0 ? 2'h0 : lvtReg_419; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_420 = 10'h1a4 == io_wrAddr_0 ? 2'h0 : lvtReg_420; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_421 = 10'h1a5 == io_wrAddr_0 ? 2'h0 : lvtReg_421; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_422 = 10'h1a6 == io_wrAddr_0 ? 2'h0 : lvtReg_422; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_423 = 10'h1a7 == io_wrAddr_0 ? 2'h0 : lvtReg_423; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_424 = 10'h1a8 == io_wrAddr_0 ? 2'h0 : lvtReg_424; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_425 = 10'h1a9 == io_wrAddr_0 ? 2'h0 : lvtReg_425; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_426 = 10'h1aa == io_wrAddr_0 ? 2'h0 : lvtReg_426; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_427 = 10'h1ab == io_wrAddr_0 ? 2'h0 : lvtReg_427; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_428 = 10'h1ac == io_wrAddr_0 ? 2'h0 : lvtReg_428; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_429 = 10'h1ad == io_wrAddr_0 ? 2'h0 : lvtReg_429; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_430 = 10'h1ae == io_wrAddr_0 ? 2'h0 : lvtReg_430; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_431 = 10'h1af == io_wrAddr_0 ? 2'h0 : lvtReg_431; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_432 = 10'h1b0 == io_wrAddr_0 ? 2'h0 : lvtReg_432; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_433 = 10'h1b1 == io_wrAddr_0 ? 2'h0 : lvtReg_433; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_434 = 10'h1b2 == io_wrAddr_0 ? 2'h0 : lvtReg_434; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_435 = 10'h1b3 == io_wrAddr_0 ? 2'h0 : lvtReg_435; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_436 = 10'h1b4 == io_wrAddr_0 ? 2'h0 : lvtReg_436; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_437 = 10'h1b5 == io_wrAddr_0 ? 2'h0 : lvtReg_437; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_438 = 10'h1b6 == io_wrAddr_0 ? 2'h0 : lvtReg_438; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_439 = 10'h1b7 == io_wrAddr_0 ? 2'h0 : lvtReg_439; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_440 = 10'h1b8 == io_wrAddr_0 ? 2'h0 : lvtReg_440; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_441 = 10'h1b9 == io_wrAddr_0 ? 2'h0 : lvtReg_441; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_442 = 10'h1ba == io_wrAddr_0 ? 2'h0 : lvtReg_442; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_443 = 10'h1bb == io_wrAddr_0 ? 2'h0 : lvtReg_443; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_444 = 10'h1bc == io_wrAddr_0 ? 2'h0 : lvtReg_444; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_445 = 10'h1bd == io_wrAddr_0 ? 2'h0 : lvtReg_445; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_446 = 10'h1be == io_wrAddr_0 ? 2'h0 : lvtReg_446; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_447 = 10'h1bf == io_wrAddr_0 ? 2'h0 : lvtReg_447; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_448 = 10'h1c0 == io_wrAddr_0 ? 2'h0 : lvtReg_448; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_449 = 10'h1c1 == io_wrAddr_0 ? 2'h0 : lvtReg_449; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_450 = 10'h1c2 == io_wrAddr_0 ? 2'h0 : lvtReg_450; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_451 = 10'h1c3 == io_wrAddr_0 ? 2'h0 : lvtReg_451; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_452 = 10'h1c4 == io_wrAddr_0 ? 2'h0 : lvtReg_452; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_453 = 10'h1c5 == io_wrAddr_0 ? 2'h0 : lvtReg_453; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_454 = 10'h1c6 == io_wrAddr_0 ? 2'h0 : lvtReg_454; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_455 = 10'h1c7 == io_wrAddr_0 ? 2'h0 : lvtReg_455; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_456 = 10'h1c8 == io_wrAddr_0 ? 2'h0 : lvtReg_456; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_457 = 10'h1c9 == io_wrAddr_0 ? 2'h0 : lvtReg_457; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_458 = 10'h1ca == io_wrAddr_0 ? 2'h0 : lvtReg_458; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_459 = 10'h1cb == io_wrAddr_0 ? 2'h0 : lvtReg_459; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_460 = 10'h1cc == io_wrAddr_0 ? 2'h0 : lvtReg_460; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_461 = 10'h1cd == io_wrAddr_0 ? 2'h0 : lvtReg_461; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_462 = 10'h1ce == io_wrAddr_0 ? 2'h0 : lvtReg_462; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_463 = 10'h1cf == io_wrAddr_0 ? 2'h0 : lvtReg_463; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_464 = 10'h1d0 == io_wrAddr_0 ? 2'h0 : lvtReg_464; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_465 = 10'h1d1 == io_wrAddr_0 ? 2'h0 : lvtReg_465; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_466 = 10'h1d2 == io_wrAddr_0 ? 2'h0 : lvtReg_466; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_467 = 10'h1d3 == io_wrAddr_0 ? 2'h0 : lvtReg_467; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_468 = 10'h1d4 == io_wrAddr_0 ? 2'h0 : lvtReg_468; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_469 = 10'h1d5 == io_wrAddr_0 ? 2'h0 : lvtReg_469; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_470 = 10'h1d6 == io_wrAddr_0 ? 2'h0 : lvtReg_470; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_471 = 10'h1d7 == io_wrAddr_0 ? 2'h0 : lvtReg_471; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_472 = 10'h1d8 == io_wrAddr_0 ? 2'h0 : lvtReg_472; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_473 = 10'h1d9 == io_wrAddr_0 ? 2'h0 : lvtReg_473; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_474 = 10'h1da == io_wrAddr_0 ? 2'h0 : lvtReg_474; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_475 = 10'h1db == io_wrAddr_0 ? 2'h0 : lvtReg_475; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_476 = 10'h1dc == io_wrAddr_0 ? 2'h0 : lvtReg_476; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_477 = 10'h1dd == io_wrAddr_0 ? 2'h0 : lvtReg_477; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_478 = 10'h1de == io_wrAddr_0 ? 2'h0 : lvtReg_478; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_479 = 10'h1df == io_wrAddr_0 ? 2'h0 : lvtReg_479; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_480 = 10'h1e0 == io_wrAddr_0 ? 2'h0 : lvtReg_480; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_481 = 10'h1e1 == io_wrAddr_0 ? 2'h0 : lvtReg_481; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_482 = 10'h1e2 == io_wrAddr_0 ? 2'h0 : lvtReg_482; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_483 = 10'h1e3 == io_wrAddr_0 ? 2'h0 : lvtReg_483; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_484 = 10'h1e4 == io_wrAddr_0 ? 2'h0 : lvtReg_484; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_485 = 10'h1e5 == io_wrAddr_0 ? 2'h0 : lvtReg_485; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_486 = 10'h1e6 == io_wrAddr_0 ? 2'h0 : lvtReg_486; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_487 = 10'h1e7 == io_wrAddr_0 ? 2'h0 : lvtReg_487; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_488 = 10'h1e8 == io_wrAddr_0 ? 2'h0 : lvtReg_488; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_489 = 10'h1e9 == io_wrAddr_0 ? 2'h0 : lvtReg_489; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_490 = 10'h1ea == io_wrAddr_0 ? 2'h0 : lvtReg_490; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_491 = 10'h1eb == io_wrAddr_0 ? 2'h0 : lvtReg_491; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_492 = 10'h1ec == io_wrAddr_0 ? 2'h0 : lvtReg_492; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_493 = 10'h1ed == io_wrAddr_0 ? 2'h0 : lvtReg_493; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_494 = 10'h1ee == io_wrAddr_0 ? 2'h0 : lvtReg_494; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_495 = 10'h1ef == io_wrAddr_0 ? 2'h0 : lvtReg_495; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_496 = 10'h1f0 == io_wrAddr_0 ? 2'h0 : lvtReg_496; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_497 = 10'h1f1 == io_wrAddr_0 ? 2'h0 : lvtReg_497; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_498 = 10'h1f2 == io_wrAddr_0 ? 2'h0 : lvtReg_498; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_499 = 10'h1f3 == io_wrAddr_0 ? 2'h0 : lvtReg_499; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_500 = 10'h1f4 == io_wrAddr_0 ? 2'h0 : lvtReg_500; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_501 = 10'h1f5 == io_wrAddr_0 ? 2'h0 : lvtReg_501; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_502 = 10'h1f6 == io_wrAddr_0 ? 2'h0 : lvtReg_502; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_503 = 10'h1f7 == io_wrAddr_0 ? 2'h0 : lvtReg_503; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_504 = 10'h1f8 == io_wrAddr_0 ? 2'h0 : lvtReg_504; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_505 = 10'h1f9 == io_wrAddr_0 ? 2'h0 : lvtReg_505; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_506 = 10'h1fa == io_wrAddr_0 ? 2'h0 : lvtReg_506; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_507 = 10'h1fb == io_wrAddr_0 ? 2'h0 : lvtReg_507; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_508 = 10'h1fc == io_wrAddr_0 ? 2'h0 : lvtReg_508; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_509 = 10'h1fd == io_wrAddr_0 ? 2'h0 : lvtReg_509; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_510 = 10'h1fe == io_wrAddr_0 ? 2'h0 : lvtReg_510; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_511 = 10'h1ff == io_wrAddr_0 ? 2'h0 : lvtReg_511; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_512 = 10'h200 == io_wrAddr_0 ? 2'h0 : lvtReg_512; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_513 = 10'h201 == io_wrAddr_0 ? 2'h0 : lvtReg_513; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_514 = 10'h202 == io_wrAddr_0 ? 2'h0 : lvtReg_514; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_515 = 10'h203 == io_wrAddr_0 ? 2'h0 : lvtReg_515; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_516 = 10'h204 == io_wrAddr_0 ? 2'h0 : lvtReg_516; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_517 = 10'h205 == io_wrAddr_0 ? 2'h0 : lvtReg_517; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_518 = 10'h206 == io_wrAddr_0 ? 2'h0 : lvtReg_518; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_519 = 10'h207 == io_wrAddr_0 ? 2'h0 : lvtReg_519; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_520 = 10'h208 == io_wrAddr_0 ? 2'h0 : lvtReg_520; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_521 = 10'h209 == io_wrAddr_0 ? 2'h0 : lvtReg_521; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_522 = 10'h20a == io_wrAddr_0 ? 2'h0 : lvtReg_522; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_523 = 10'h20b == io_wrAddr_0 ? 2'h0 : lvtReg_523; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_524 = 10'h20c == io_wrAddr_0 ? 2'h0 : lvtReg_524; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_525 = 10'h20d == io_wrAddr_0 ? 2'h0 : lvtReg_525; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_526 = 10'h20e == io_wrAddr_0 ? 2'h0 : lvtReg_526; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_527 = 10'h20f == io_wrAddr_0 ? 2'h0 : lvtReg_527; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_528 = 10'h210 == io_wrAddr_0 ? 2'h0 : lvtReg_528; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_529 = 10'h211 == io_wrAddr_0 ? 2'h0 : lvtReg_529; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_530 = 10'h212 == io_wrAddr_0 ? 2'h0 : lvtReg_530; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_531 = 10'h213 == io_wrAddr_0 ? 2'h0 : lvtReg_531; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_532 = 10'h214 == io_wrAddr_0 ? 2'h0 : lvtReg_532; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_533 = 10'h215 == io_wrAddr_0 ? 2'h0 : lvtReg_533; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_534 = 10'h216 == io_wrAddr_0 ? 2'h0 : lvtReg_534; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_535 = 10'h217 == io_wrAddr_0 ? 2'h0 : lvtReg_535; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_536 = 10'h218 == io_wrAddr_0 ? 2'h0 : lvtReg_536; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_537 = 10'h219 == io_wrAddr_0 ? 2'h0 : lvtReg_537; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_538 = 10'h21a == io_wrAddr_0 ? 2'h0 : lvtReg_538; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_539 = 10'h21b == io_wrAddr_0 ? 2'h0 : lvtReg_539; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_540 = 10'h21c == io_wrAddr_0 ? 2'h0 : lvtReg_540; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_541 = 10'h21d == io_wrAddr_0 ? 2'h0 : lvtReg_541; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_542 = 10'h21e == io_wrAddr_0 ? 2'h0 : lvtReg_542; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_543 = 10'h21f == io_wrAddr_0 ? 2'h0 : lvtReg_543; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_544 = 10'h220 == io_wrAddr_0 ? 2'h0 : lvtReg_544; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_545 = 10'h221 == io_wrAddr_0 ? 2'h0 : lvtReg_545; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_546 = 10'h222 == io_wrAddr_0 ? 2'h0 : lvtReg_546; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_547 = 10'h223 == io_wrAddr_0 ? 2'h0 : lvtReg_547; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_548 = 10'h224 == io_wrAddr_0 ? 2'h0 : lvtReg_548; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_549 = 10'h225 == io_wrAddr_0 ? 2'h0 : lvtReg_549; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_550 = 10'h226 == io_wrAddr_0 ? 2'h0 : lvtReg_550; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_551 = 10'h227 == io_wrAddr_0 ? 2'h0 : lvtReg_551; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_552 = 10'h228 == io_wrAddr_0 ? 2'h0 : lvtReg_552; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_553 = 10'h229 == io_wrAddr_0 ? 2'h0 : lvtReg_553; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_554 = 10'h22a == io_wrAddr_0 ? 2'h0 : lvtReg_554; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_555 = 10'h22b == io_wrAddr_0 ? 2'h0 : lvtReg_555; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_556 = 10'h22c == io_wrAddr_0 ? 2'h0 : lvtReg_556; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_557 = 10'h22d == io_wrAddr_0 ? 2'h0 : lvtReg_557; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_558 = 10'h22e == io_wrAddr_0 ? 2'h0 : lvtReg_558; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_559 = 10'h22f == io_wrAddr_0 ? 2'h0 : lvtReg_559; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_560 = 10'h230 == io_wrAddr_0 ? 2'h0 : lvtReg_560; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_561 = 10'h231 == io_wrAddr_0 ? 2'h0 : lvtReg_561; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_562 = 10'h232 == io_wrAddr_0 ? 2'h0 : lvtReg_562; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_563 = 10'h233 == io_wrAddr_0 ? 2'h0 : lvtReg_563; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_564 = 10'h234 == io_wrAddr_0 ? 2'h0 : lvtReg_564; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_565 = 10'h235 == io_wrAddr_0 ? 2'h0 : lvtReg_565; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_566 = 10'h236 == io_wrAddr_0 ? 2'h0 : lvtReg_566; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_567 = 10'h237 == io_wrAddr_0 ? 2'h0 : lvtReg_567; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_568 = 10'h238 == io_wrAddr_0 ? 2'h0 : lvtReg_568; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_569 = 10'h239 == io_wrAddr_0 ? 2'h0 : lvtReg_569; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_570 = 10'h23a == io_wrAddr_0 ? 2'h0 : lvtReg_570; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_571 = 10'h23b == io_wrAddr_0 ? 2'h0 : lvtReg_571; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_572 = 10'h23c == io_wrAddr_0 ? 2'h0 : lvtReg_572; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_573 = 10'h23d == io_wrAddr_0 ? 2'h0 : lvtReg_573; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_574 = 10'h23e == io_wrAddr_0 ? 2'h0 : lvtReg_574; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_575 = 10'h23f == io_wrAddr_0 ? 2'h0 : lvtReg_575; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_576 = 10'h240 == io_wrAddr_0 ? 2'h0 : lvtReg_576; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_577 = 10'h241 == io_wrAddr_0 ? 2'h0 : lvtReg_577; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_578 = 10'h242 == io_wrAddr_0 ? 2'h0 : lvtReg_578; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_579 = 10'h243 == io_wrAddr_0 ? 2'h0 : lvtReg_579; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_580 = 10'h244 == io_wrAddr_0 ? 2'h0 : lvtReg_580; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_581 = 10'h245 == io_wrAddr_0 ? 2'h0 : lvtReg_581; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_582 = 10'h246 == io_wrAddr_0 ? 2'h0 : lvtReg_582; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_583 = 10'h247 == io_wrAddr_0 ? 2'h0 : lvtReg_583; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_584 = 10'h248 == io_wrAddr_0 ? 2'h0 : lvtReg_584; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_585 = 10'h249 == io_wrAddr_0 ? 2'h0 : lvtReg_585; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_586 = 10'h24a == io_wrAddr_0 ? 2'h0 : lvtReg_586; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_587 = 10'h24b == io_wrAddr_0 ? 2'h0 : lvtReg_587; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_588 = 10'h24c == io_wrAddr_0 ? 2'h0 : lvtReg_588; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_589 = 10'h24d == io_wrAddr_0 ? 2'h0 : lvtReg_589; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_590 = 10'h24e == io_wrAddr_0 ? 2'h0 : lvtReg_590; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_591 = 10'h24f == io_wrAddr_0 ? 2'h0 : lvtReg_591; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_592 = 10'h250 == io_wrAddr_0 ? 2'h0 : lvtReg_592; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_593 = 10'h251 == io_wrAddr_0 ? 2'h0 : lvtReg_593; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_594 = 10'h252 == io_wrAddr_0 ? 2'h0 : lvtReg_594; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_595 = 10'h253 == io_wrAddr_0 ? 2'h0 : lvtReg_595; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_596 = 10'h254 == io_wrAddr_0 ? 2'h0 : lvtReg_596; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_597 = 10'h255 == io_wrAddr_0 ? 2'h0 : lvtReg_597; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_598 = 10'h256 == io_wrAddr_0 ? 2'h0 : lvtReg_598; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_599 = 10'h257 == io_wrAddr_0 ? 2'h0 : lvtReg_599; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_600 = 10'h258 == io_wrAddr_0 ? 2'h0 : lvtReg_600; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_601 = 10'h259 == io_wrAddr_0 ? 2'h0 : lvtReg_601; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_602 = 10'h25a == io_wrAddr_0 ? 2'h0 : lvtReg_602; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_603 = 10'h25b == io_wrAddr_0 ? 2'h0 : lvtReg_603; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_604 = 10'h25c == io_wrAddr_0 ? 2'h0 : lvtReg_604; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_605 = 10'h25d == io_wrAddr_0 ? 2'h0 : lvtReg_605; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_606 = 10'h25e == io_wrAddr_0 ? 2'h0 : lvtReg_606; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_607 = 10'h25f == io_wrAddr_0 ? 2'h0 : lvtReg_607; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_608 = 10'h260 == io_wrAddr_0 ? 2'h0 : lvtReg_608; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_609 = 10'h261 == io_wrAddr_0 ? 2'h0 : lvtReg_609; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_610 = 10'h262 == io_wrAddr_0 ? 2'h0 : lvtReg_610; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_611 = 10'h263 == io_wrAddr_0 ? 2'h0 : lvtReg_611; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_612 = 10'h264 == io_wrAddr_0 ? 2'h0 : lvtReg_612; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_613 = 10'h265 == io_wrAddr_0 ? 2'h0 : lvtReg_613; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_614 = 10'h266 == io_wrAddr_0 ? 2'h0 : lvtReg_614; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_615 = 10'h267 == io_wrAddr_0 ? 2'h0 : lvtReg_615; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_616 = 10'h268 == io_wrAddr_0 ? 2'h0 : lvtReg_616; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_617 = 10'h269 == io_wrAddr_0 ? 2'h0 : lvtReg_617; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_618 = 10'h26a == io_wrAddr_0 ? 2'h0 : lvtReg_618; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_619 = 10'h26b == io_wrAddr_0 ? 2'h0 : lvtReg_619; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_620 = 10'h26c == io_wrAddr_0 ? 2'h0 : lvtReg_620; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_621 = 10'h26d == io_wrAddr_0 ? 2'h0 : lvtReg_621; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_622 = 10'h26e == io_wrAddr_0 ? 2'h0 : lvtReg_622; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_623 = 10'h26f == io_wrAddr_0 ? 2'h0 : lvtReg_623; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_624 = 10'h270 == io_wrAddr_0 ? 2'h0 : lvtReg_624; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_625 = 10'h271 == io_wrAddr_0 ? 2'h0 : lvtReg_625; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_626 = 10'h272 == io_wrAddr_0 ? 2'h0 : lvtReg_626; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_627 = 10'h273 == io_wrAddr_0 ? 2'h0 : lvtReg_627; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_628 = 10'h274 == io_wrAddr_0 ? 2'h0 : lvtReg_628; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_629 = 10'h275 == io_wrAddr_0 ? 2'h0 : lvtReg_629; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_630 = 10'h276 == io_wrAddr_0 ? 2'h0 : lvtReg_630; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_631 = 10'h277 == io_wrAddr_0 ? 2'h0 : lvtReg_631; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_632 = 10'h278 == io_wrAddr_0 ? 2'h0 : lvtReg_632; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_633 = 10'h279 == io_wrAddr_0 ? 2'h0 : lvtReg_633; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_634 = 10'h27a == io_wrAddr_0 ? 2'h0 : lvtReg_634; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_635 = 10'h27b == io_wrAddr_0 ? 2'h0 : lvtReg_635; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_636 = 10'h27c == io_wrAddr_0 ? 2'h0 : lvtReg_636; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_637 = 10'h27d == io_wrAddr_0 ? 2'h0 : lvtReg_637; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_638 = 10'h27e == io_wrAddr_0 ? 2'h0 : lvtReg_638; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_639 = 10'h27f == io_wrAddr_0 ? 2'h0 : lvtReg_639; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_640 = 10'h280 == io_wrAddr_0 ? 2'h0 : lvtReg_640; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_641 = 10'h281 == io_wrAddr_0 ? 2'h0 : lvtReg_641; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_642 = 10'h282 == io_wrAddr_0 ? 2'h0 : lvtReg_642; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_643 = 10'h283 == io_wrAddr_0 ? 2'h0 : lvtReg_643; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_644 = 10'h284 == io_wrAddr_0 ? 2'h0 : lvtReg_644; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_645 = 10'h285 == io_wrAddr_0 ? 2'h0 : lvtReg_645; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_646 = 10'h286 == io_wrAddr_0 ? 2'h0 : lvtReg_646; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_647 = 10'h287 == io_wrAddr_0 ? 2'h0 : lvtReg_647; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_648 = 10'h288 == io_wrAddr_0 ? 2'h0 : lvtReg_648; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_649 = 10'h289 == io_wrAddr_0 ? 2'h0 : lvtReg_649; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_650 = 10'h28a == io_wrAddr_0 ? 2'h0 : lvtReg_650; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_651 = 10'h28b == io_wrAddr_0 ? 2'h0 : lvtReg_651; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_652 = 10'h28c == io_wrAddr_0 ? 2'h0 : lvtReg_652; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_653 = 10'h28d == io_wrAddr_0 ? 2'h0 : lvtReg_653; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_654 = 10'h28e == io_wrAddr_0 ? 2'h0 : lvtReg_654; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_655 = 10'h28f == io_wrAddr_0 ? 2'h0 : lvtReg_655; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_656 = 10'h290 == io_wrAddr_0 ? 2'h0 : lvtReg_656; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_657 = 10'h291 == io_wrAddr_0 ? 2'h0 : lvtReg_657; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_658 = 10'h292 == io_wrAddr_0 ? 2'h0 : lvtReg_658; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_659 = 10'h293 == io_wrAddr_0 ? 2'h0 : lvtReg_659; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_660 = 10'h294 == io_wrAddr_0 ? 2'h0 : lvtReg_660; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_661 = 10'h295 == io_wrAddr_0 ? 2'h0 : lvtReg_661; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_662 = 10'h296 == io_wrAddr_0 ? 2'h0 : lvtReg_662; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_663 = 10'h297 == io_wrAddr_0 ? 2'h0 : lvtReg_663; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_664 = 10'h298 == io_wrAddr_0 ? 2'h0 : lvtReg_664; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_665 = 10'h299 == io_wrAddr_0 ? 2'h0 : lvtReg_665; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_666 = 10'h29a == io_wrAddr_0 ? 2'h0 : lvtReg_666; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_667 = 10'h29b == io_wrAddr_0 ? 2'h0 : lvtReg_667; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_668 = 10'h29c == io_wrAddr_0 ? 2'h0 : lvtReg_668; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_669 = 10'h29d == io_wrAddr_0 ? 2'h0 : lvtReg_669; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_670 = 10'h29e == io_wrAddr_0 ? 2'h0 : lvtReg_670; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_671 = 10'h29f == io_wrAddr_0 ? 2'h0 : lvtReg_671; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_672 = 10'h2a0 == io_wrAddr_0 ? 2'h0 : lvtReg_672; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_673 = 10'h2a1 == io_wrAddr_0 ? 2'h0 : lvtReg_673; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_674 = 10'h2a2 == io_wrAddr_0 ? 2'h0 : lvtReg_674; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_675 = 10'h2a3 == io_wrAddr_0 ? 2'h0 : lvtReg_675; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_676 = 10'h2a4 == io_wrAddr_0 ? 2'h0 : lvtReg_676; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_677 = 10'h2a5 == io_wrAddr_0 ? 2'h0 : lvtReg_677; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_678 = 10'h2a6 == io_wrAddr_0 ? 2'h0 : lvtReg_678; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_679 = 10'h2a7 == io_wrAddr_0 ? 2'h0 : lvtReg_679; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_680 = 10'h2a8 == io_wrAddr_0 ? 2'h0 : lvtReg_680; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_681 = 10'h2a9 == io_wrAddr_0 ? 2'h0 : lvtReg_681; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_682 = 10'h2aa == io_wrAddr_0 ? 2'h0 : lvtReg_682; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_683 = 10'h2ab == io_wrAddr_0 ? 2'h0 : lvtReg_683; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_684 = 10'h2ac == io_wrAddr_0 ? 2'h0 : lvtReg_684; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_685 = 10'h2ad == io_wrAddr_0 ? 2'h0 : lvtReg_685; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_686 = 10'h2ae == io_wrAddr_0 ? 2'h0 : lvtReg_686; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_687 = 10'h2af == io_wrAddr_0 ? 2'h0 : lvtReg_687; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_688 = 10'h2b0 == io_wrAddr_0 ? 2'h0 : lvtReg_688; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_689 = 10'h2b1 == io_wrAddr_0 ? 2'h0 : lvtReg_689; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_690 = 10'h2b2 == io_wrAddr_0 ? 2'h0 : lvtReg_690; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_691 = 10'h2b3 == io_wrAddr_0 ? 2'h0 : lvtReg_691; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_692 = 10'h2b4 == io_wrAddr_0 ? 2'h0 : lvtReg_692; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_693 = 10'h2b5 == io_wrAddr_0 ? 2'h0 : lvtReg_693; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_694 = 10'h2b6 == io_wrAddr_0 ? 2'h0 : lvtReg_694; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_695 = 10'h2b7 == io_wrAddr_0 ? 2'h0 : lvtReg_695; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_696 = 10'h2b8 == io_wrAddr_0 ? 2'h0 : lvtReg_696; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_697 = 10'h2b9 == io_wrAddr_0 ? 2'h0 : lvtReg_697; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_698 = 10'h2ba == io_wrAddr_0 ? 2'h0 : lvtReg_698; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_699 = 10'h2bb == io_wrAddr_0 ? 2'h0 : lvtReg_699; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_700 = 10'h2bc == io_wrAddr_0 ? 2'h0 : lvtReg_700; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_701 = 10'h2bd == io_wrAddr_0 ? 2'h0 : lvtReg_701; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_702 = 10'h2be == io_wrAddr_0 ? 2'h0 : lvtReg_702; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_703 = 10'h2bf == io_wrAddr_0 ? 2'h0 : lvtReg_703; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_704 = 10'h2c0 == io_wrAddr_0 ? 2'h0 : lvtReg_704; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_705 = 10'h2c1 == io_wrAddr_0 ? 2'h0 : lvtReg_705; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_706 = 10'h2c2 == io_wrAddr_0 ? 2'h0 : lvtReg_706; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_707 = 10'h2c3 == io_wrAddr_0 ? 2'h0 : lvtReg_707; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_708 = 10'h2c4 == io_wrAddr_0 ? 2'h0 : lvtReg_708; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_709 = 10'h2c5 == io_wrAddr_0 ? 2'h0 : lvtReg_709; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_710 = 10'h2c6 == io_wrAddr_0 ? 2'h0 : lvtReg_710; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_711 = 10'h2c7 == io_wrAddr_0 ? 2'h0 : lvtReg_711; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_712 = 10'h2c8 == io_wrAddr_0 ? 2'h0 : lvtReg_712; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_713 = 10'h2c9 == io_wrAddr_0 ? 2'h0 : lvtReg_713; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_714 = 10'h2ca == io_wrAddr_0 ? 2'h0 : lvtReg_714; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_715 = 10'h2cb == io_wrAddr_0 ? 2'h0 : lvtReg_715; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_716 = 10'h2cc == io_wrAddr_0 ? 2'h0 : lvtReg_716; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_717 = 10'h2cd == io_wrAddr_0 ? 2'h0 : lvtReg_717; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_718 = 10'h2ce == io_wrAddr_0 ? 2'h0 : lvtReg_718; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_719 = 10'h2cf == io_wrAddr_0 ? 2'h0 : lvtReg_719; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_720 = 10'h2d0 == io_wrAddr_0 ? 2'h0 : lvtReg_720; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_721 = 10'h2d1 == io_wrAddr_0 ? 2'h0 : lvtReg_721; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_722 = 10'h2d2 == io_wrAddr_0 ? 2'h0 : lvtReg_722; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_723 = 10'h2d3 == io_wrAddr_0 ? 2'h0 : lvtReg_723; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_724 = 10'h2d4 == io_wrAddr_0 ? 2'h0 : lvtReg_724; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_725 = 10'h2d5 == io_wrAddr_0 ? 2'h0 : lvtReg_725; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_726 = 10'h2d6 == io_wrAddr_0 ? 2'h0 : lvtReg_726; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_727 = 10'h2d7 == io_wrAddr_0 ? 2'h0 : lvtReg_727; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_728 = 10'h2d8 == io_wrAddr_0 ? 2'h0 : lvtReg_728; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_729 = 10'h2d9 == io_wrAddr_0 ? 2'h0 : lvtReg_729; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_730 = 10'h2da == io_wrAddr_0 ? 2'h0 : lvtReg_730; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_731 = 10'h2db == io_wrAddr_0 ? 2'h0 : lvtReg_731; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_732 = 10'h2dc == io_wrAddr_0 ? 2'h0 : lvtReg_732; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_733 = 10'h2dd == io_wrAddr_0 ? 2'h0 : lvtReg_733; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_734 = 10'h2de == io_wrAddr_0 ? 2'h0 : lvtReg_734; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_735 = 10'h2df == io_wrAddr_0 ? 2'h0 : lvtReg_735; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_736 = 10'h2e0 == io_wrAddr_0 ? 2'h0 : lvtReg_736; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_737 = 10'h2e1 == io_wrAddr_0 ? 2'h0 : lvtReg_737; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_738 = 10'h2e2 == io_wrAddr_0 ? 2'h0 : lvtReg_738; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_739 = 10'h2e3 == io_wrAddr_0 ? 2'h0 : lvtReg_739; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_740 = 10'h2e4 == io_wrAddr_0 ? 2'h0 : lvtReg_740; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_741 = 10'h2e5 == io_wrAddr_0 ? 2'h0 : lvtReg_741; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_742 = 10'h2e6 == io_wrAddr_0 ? 2'h0 : lvtReg_742; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_743 = 10'h2e7 == io_wrAddr_0 ? 2'h0 : lvtReg_743; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_744 = 10'h2e8 == io_wrAddr_0 ? 2'h0 : lvtReg_744; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_745 = 10'h2e9 == io_wrAddr_0 ? 2'h0 : lvtReg_745; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_746 = 10'h2ea == io_wrAddr_0 ? 2'h0 : lvtReg_746; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_747 = 10'h2eb == io_wrAddr_0 ? 2'h0 : lvtReg_747; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_748 = 10'h2ec == io_wrAddr_0 ? 2'h0 : lvtReg_748; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_749 = 10'h2ed == io_wrAddr_0 ? 2'h0 : lvtReg_749; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_750 = 10'h2ee == io_wrAddr_0 ? 2'h0 : lvtReg_750; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_751 = 10'h2ef == io_wrAddr_0 ? 2'h0 : lvtReg_751; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_752 = 10'h2f0 == io_wrAddr_0 ? 2'h0 : lvtReg_752; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_753 = 10'h2f1 == io_wrAddr_0 ? 2'h0 : lvtReg_753; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_754 = 10'h2f2 == io_wrAddr_0 ? 2'h0 : lvtReg_754; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_755 = 10'h2f3 == io_wrAddr_0 ? 2'h0 : lvtReg_755; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_756 = 10'h2f4 == io_wrAddr_0 ? 2'h0 : lvtReg_756; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_757 = 10'h2f5 == io_wrAddr_0 ? 2'h0 : lvtReg_757; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_758 = 10'h2f6 == io_wrAddr_0 ? 2'h0 : lvtReg_758; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_759 = 10'h2f7 == io_wrAddr_0 ? 2'h0 : lvtReg_759; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_760 = 10'h2f8 == io_wrAddr_0 ? 2'h0 : lvtReg_760; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_761 = 10'h2f9 == io_wrAddr_0 ? 2'h0 : lvtReg_761; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_762 = 10'h2fa == io_wrAddr_0 ? 2'h0 : lvtReg_762; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_763 = 10'h2fb == io_wrAddr_0 ? 2'h0 : lvtReg_763; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_764 = 10'h2fc == io_wrAddr_0 ? 2'h0 : lvtReg_764; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_765 = 10'h2fd == io_wrAddr_0 ? 2'h0 : lvtReg_765; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_766 = 10'h2fe == io_wrAddr_0 ? 2'h0 : lvtReg_766; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_767 = 10'h2ff == io_wrAddr_0 ? 2'h0 : lvtReg_767; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_768 = 10'h300 == io_wrAddr_0 ? 2'h0 : lvtReg_768; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_769 = 10'h301 == io_wrAddr_0 ? 2'h0 : lvtReg_769; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_770 = 10'h302 == io_wrAddr_0 ? 2'h0 : lvtReg_770; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_771 = 10'h303 == io_wrAddr_0 ? 2'h0 : lvtReg_771; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_772 = 10'h304 == io_wrAddr_0 ? 2'h0 : lvtReg_772; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_773 = 10'h305 == io_wrAddr_0 ? 2'h0 : lvtReg_773; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_774 = 10'h306 == io_wrAddr_0 ? 2'h0 : lvtReg_774; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_775 = 10'h307 == io_wrAddr_0 ? 2'h0 : lvtReg_775; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_776 = 10'h308 == io_wrAddr_0 ? 2'h0 : lvtReg_776; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_777 = 10'h309 == io_wrAddr_0 ? 2'h0 : lvtReg_777; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_778 = 10'h30a == io_wrAddr_0 ? 2'h0 : lvtReg_778; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_779 = 10'h30b == io_wrAddr_0 ? 2'h0 : lvtReg_779; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_780 = 10'h30c == io_wrAddr_0 ? 2'h0 : lvtReg_780; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_781 = 10'h30d == io_wrAddr_0 ? 2'h0 : lvtReg_781; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_782 = 10'h30e == io_wrAddr_0 ? 2'h0 : lvtReg_782; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_783 = 10'h30f == io_wrAddr_0 ? 2'h0 : lvtReg_783; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_784 = 10'h310 == io_wrAddr_0 ? 2'h0 : lvtReg_784; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_785 = 10'h311 == io_wrAddr_0 ? 2'h0 : lvtReg_785; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_786 = 10'h312 == io_wrAddr_0 ? 2'h0 : lvtReg_786; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_787 = 10'h313 == io_wrAddr_0 ? 2'h0 : lvtReg_787; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_788 = 10'h314 == io_wrAddr_0 ? 2'h0 : lvtReg_788; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_789 = 10'h315 == io_wrAddr_0 ? 2'h0 : lvtReg_789; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_790 = 10'h316 == io_wrAddr_0 ? 2'h0 : lvtReg_790; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_791 = 10'h317 == io_wrAddr_0 ? 2'h0 : lvtReg_791; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_792 = 10'h318 == io_wrAddr_0 ? 2'h0 : lvtReg_792; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_793 = 10'h319 == io_wrAddr_0 ? 2'h0 : lvtReg_793; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_794 = 10'h31a == io_wrAddr_0 ? 2'h0 : lvtReg_794; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_795 = 10'h31b == io_wrAddr_0 ? 2'h0 : lvtReg_795; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_796 = 10'h31c == io_wrAddr_0 ? 2'h0 : lvtReg_796; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_797 = 10'h31d == io_wrAddr_0 ? 2'h0 : lvtReg_797; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_798 = 10'h31e == io_wrAddr_0 ? 2'h0 : lvtReg_798; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_799 = 10'h31f == io_wrAddr_0 ? 2'h0 : lvtReg_799; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_800 = 10'h320 == io_wrAddr_0 ? 2'h0 : lvtReg_800; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_801 = 10'h321 == io_wrAddr_0 ? 2'h0 : lvtReg_801; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_802 = 10'h322 == io_wrAddr_0 ? 2'h0 : lvtReg_802; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_803 = 10'h323 == io_wrAddr_0 ? 2'h0 : lvtReg_803; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_804 = 10'h324 == io_wrAddr_0 ? 2'h0 : lvtReg_804; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_805 = 10'h325 == io_wrAddr_0 ? 2'h0 : lvtReg_805; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_806 = 10'h326 == io_wrAddr_0 ? 2'h0 : lvtReg_806; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_807 = 10'h327 == io_wrAddr_0 ? 2'h0 : lvtReg_807; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_808 = 10'h328 == io_wrAddr_0 ? 2'h0 : lvtReg_808; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_809 = 10'h329 == io_wrAddr_0 ? 2'h0 : lvtReg_809; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_810 = 10'h32a == io_wrAddr_0 ? 2'h0 : lvtReg_810; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_811 = 10'h32b == io_wrAddr_0 ? 2'h0 : lvtReg_811; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_812 = 10'h32c == io_wrAddr_0 ? 2'h0 : lvtReg_812; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_813 = 10'h32d == io_wrAddr_0 ? 2'h0 : lvtReg_813; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_814 = 10'h32e == io_wrAddr_0 ? 2'h0 : lvtReg_814; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_815 = 10'h32f == io_wrAddr_0 ? 2'h0 : lvtReg_815; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_816 = 10'h330 == io_wrAddr_0 ? 2'h0 : lvtReg_816; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_817 = 10'h331 == io_wrAddr_0 ? 2'h0 : lvtReg_817; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_818 = 10'h332 == io_wrAddr_0 ? 2'h0 : lvtReg_818; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_819 = 10'h333 == io_wrAddr_0 ? 2'h0 : lvtReg_819; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_820 = 10'h334 == io_wrAddr_0 ? 2'h0 : lvtReg_820; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_821 = 10'h335 == io_wrAddr_0 ? 2'h0 : lvtReg_821; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_822 = 10'h336 == io_wrAddr_0 ? 2'h0 : lvtReg_822; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_823 = 10'h337 == io_wrAddr_0 ? 2'h0 : lvtReg_823; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_824 = 10'h338 == io_wrAddr_0 ? 2'h0 : lvtReg_824; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_825 = 10'h339 == io_wrAddr_0 ? 2'h0 : lvtReg_825; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_826 = 10'h33a == io_wrAddr_0 ? 2'h0 : lvtReg_826; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_827 = 10'h33b == io_wrAddr_0 ? 2'h0 : lvtReg_827; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_828 = 10'h33c == io_wrAddr_0 ? 2'h0 : lvtReg_828; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_829 = 10'h33d == io_wrAddr_0 ? 2'h0 : lvtReg_829; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_830 = 10'h33e == io_wrAddr_0 ? 2'h0 : lvtReg_830; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_831 = 10'h33f == io_wrAddr_0 ? 2'h0 : lvtReg_831; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_832 = 10'h340 == io_wrAddr_0 ? 2'h0 : lvtReg_832; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_833 = 10'h341 == io_wrAddr_0 ? 2'h0 : lvtReg_833; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_834 = 10'h342 == io_wrAddr_0 ? 2'h0 : lvtReg_834; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_835 = 10'h343 == io_wrAddr_0 ? 2'h0 : lvtReg_835; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_836 = 10'h344 == io_wrAddr_0 ? 2'h0 : lvtReg_836; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_837 = 10'h345 == io_wrAddr_0 ? 2'h0 : lvtReg_837; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_838 = 10'h346 == io_wrAddr_0 ? 2'h0 : lvtReg_838; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_839 = 10'h347 == io_wrAddr_0 ? 2'h0 : lvtReg_839; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_840 = 10'h348 == io_wrAddr_0 ? 2'h0 : lvtReg_840; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_841 = 10'h349 == io_wrAddr_0 ? 2'h0 : lvtReg_841; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_842 = 10'h34a == io_wrAddr_0 ? 2'h0 : lvtReg_842; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_843 = 10'h34b == io_wrAddr_0 ? 2'h0 : lvtReg_843; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_844 = 10'h34c == io_wrAddr_0 ? 2'h0 : lvtReg_844; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_845 = 10'h34d == io_wrAddr_0 ? 2'h0 : lvtReg_845; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_846 = 10'h34e == io_wrAddr_0 ? 2'h0 : lvtReg_846; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_847 = 10'h34f == io_wrAddr_0 ? 2'h0 : lvtReg_847; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_848 = 10'h350 == io_wrAddr_0 ? 2'h0 : lvtReg_848; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_849 = 10'h351 == io_wrAddr_0 ? 2'h0 : lvtReg_849; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_850 = 10'h352 == io_wrAddr_0 ? 2'h0 : lvtReg_850; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_851 = 10'h353 == io_wrAddr_0 ? 2'h0 : lvtReg_851; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_852 = 10'h354 == io_wrAddr_0 ? 2'h0 : lvtReg_852; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_853 = 10'h355 == io_wrAddr_0 ? 2'h0 : lvtReg_853; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_854 = 10'h356 == io_wrAddr_0 ? 2'h0 : lvtReg_854; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_855 = 10'h357 == io_wrAddr_0 ? 2'h0 : lvtReg_855; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_856 = 10'h358 == io_wrAddr_0 ? 2'h0 : lvtReg_856; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_857 = 10'h359 == io_wrAddr_0 ? 2'h0 : lvtReg_857; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_858 = 10'h35a == io_wrAddr_0 ? 2'h0 : lvtReg_858; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_859 = 10'h35b == io_wrAddr_0 ? 2'h0 : lvtReg_859; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_860 = 10'h35c == io_wrAddr_0 ? 2'h0 : lvtReg_860; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_861 = 10'h35d == io_wrAddr_0 ? 2'h0 : lvtReg_861; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_862 = 10'h35e == io_wrAddr_0 ? 2'h0 : lvtReg_862; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_863 = 10'h35f == io_wrAddr_0 ? 2'h0 : lvtReg_863; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_864 = 10'h360 == io_wrAddr_0 ? 2'h0 : lvtReg_864; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_865 = 10'h361 == io_wrAddr_0 ? 2'h0 : lvtReg_865; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_866 = 10'h362 == io_wrAddr_0 ? 2'h0 : lvtReg_866; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_867 = 10'h363 == io_wrAddr_0 ? 2'h0 : lvtReg_867; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_868 = 10'h364 == io_wrAddr_0 ? 2'h0 : lvtReg_868; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_869 = 10'h365 == io_wrAddr_0 ? 2'h0 : lvtReg_869; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_870 = 10'h366 == io_wrAddr_0 ? 2'h0 : lvtReg_870; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_871 = 10'h367 == io_wrAddr_0 ? 2'h0 : lvtReg_871; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_872 = 10'h368 == io_wrAddr_0 ? 2'h0 : lvtReg_872; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_873 = 10'h369 == io_wrAddr_0 ? 2'h0 : lvtReg_873; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_874 = 10'h36a == io_wrAddr_0 ? 2'h0 : lvtReg_874; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_875 = 10'h36b == io_wrAddr_0 ? 2'h0 : lvtReg_875; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_876 = 10'h36c == io_wrAddr_0 ? 2'h0 : lvtReg_876; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_877 = 10'h36d == io_wrAddr_0 ? 2'h0 : lvtReg_877; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_878 = 10'h36e == io_wrAddr_0 ? 2'h0 : lvtReg_878; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_879 = 10'h36f == io_wrAddr_0 ? 2'h0 : lvtReg_879; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_880 = 10'h370 == io_wrAddr_0 ? 2'h0 : lvtReg_880; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_881 = 10'h371 == io_wrAddr_0 ? 2'h0 : lvtReg_881; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_882 = 10'h372 == io_wrAddr_0 ? 2'h0 : lvtReg_882; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_883 = 10'h373 == io_wrAddr_0 ? 2'h0 : lvtReg_883; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_884 = 10'h374 == io_wrAddr_0 ? 2'h0 : lvtReg_884; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_885 = 10'h375 == io_wrAddr_0 ? 2'h0 : lvtReg_885; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_886 = 10'h376 == io_wrAddr_0 ? 2'h0 : lvtReg_886; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_887 = 10'h377 == io_wrAddr_0 ? 2'h0 : lvtReg_887; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_888 = 10'h378 == io_wrAddr_0 ? 2'h0 : lvtReg_888; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_889 = 10'h379 == io_wrAddr_0 ? 2'h0 : lvtReg_889; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_890 = 10'h37a == io_wrAddr_0 ? 2'h0 : lvtReg_890; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_891 = 10'h37b == io_wrAddr_0 ? 2'h0 : lvtReg_891; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_892 = 10'h37c == io_wrAddr_0 ? 2'h0 : lvtReg_892; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_893 = 10'h37d == io_wrAddr_0 ? 2'h0 : lvtReg_893; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_894 = 10'h37e == io_wrAddr_0 ? 2'h0 : lvtReg_894; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_895 = 10'h37f == io_wrAddr_0 ? 2'h0 : lvtReg_895; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_896 = 10'h380 == io_wrAddr_0 ? 2'h0 : lvtReg_896; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_897 = 10'h381 == io_wrAddr_0 ? 2'h0 : lvtReg_897; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_898 = 10'h382 == io_wrAddr_0 ? 2'h0 : lvtReg_898; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_899 = 10'h383 == io_wrAddr_0 ? 2'h0 : lvtReg_899; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_900 = 10'h384 == io_wrAddr_0 ? 2'h0 : lvtReg_900; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_901 = 10'h385 == io_wrAddr_0 ? 2'h0 : lvtReg_901; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_902 = 10'h386 == io_wrAddr_0 ? 2'h0 : lvtReg_902; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_903 = 10'h387 == io_wrAddr_0 ? 2'h0 : lvtReg_903; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_904 = 10'h388 == io_wrAddr_0 ? 2'h0 : lvtReg_904; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_905 = 10'h389 == io_wrAddr_0 ? 2'h0 : lvtReg_905; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_906 = 10'h38a == io_wrAddr_0 ? 2'h0 : lvtReg_906; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_907 = 10'h38b == io_wrAddr_0 ? 2'h0 : lvtReg_907; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_908 = 10'h38c == io_wrAddr_0 ? 2'h0 : lvtReg_908; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_909 = 10'h38d == io_wrAddr_0 ? 2'h0 : lvtReg_909; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_910 = 10'h38e == io_wrAddr_0 ? 2'h0 : lvtReg_910; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_911 = 10'h38f == io_wrAddr_0 ? 2'h0 : lvtReg_911; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_912 = 10'h390 == io_wrAddr_0 ? 2'h0 : lvtReg_912; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_913 = 10'h391 == io_wrAddr_0 ? 2'h0 : lvtReg_913; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_914 = 10'h392 == io_wrAddr_0 ? 2'h0 : lvtReg_914; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_915 = 10'h393 == io_wrAddr_0 ? 2'h0 : lvtReg_915; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_916 = 10'h394 == io_wrAddr_0 ? 2'h0 : lvtReg_916; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_917 = 10'h395 == io_wrAddr_0 ? 2'h0 : lvtReg_917; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_918 = 10'h396 == io_wrAddr_0 ? 2'h0 : lvtReg_918; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_919 = 10'h397 == io_wrAddr_0 ? 2'h0 : lvtReg_919; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_920 = 10'h398 == io_wrAddr_0 ? 2'h0 : lvtReg_920; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_921 = 10'h399 == io_wrAddr_0 ? 2'h0 : lvtReg_921; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_922 = 10'h39a == io_wrAddr_0 ? 2'h0 : lvtReg_922; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_923 = 10'h39b == io_wrAddr_0 ? 2'h0 : lvtReg_923; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_924 = 10'h39c == io_wrAddr_0 ? 2'h0 : lvtReg_924; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_925 = 10'h39d == io_wrAddr_0 ? 2'h0 : lvtReg_925; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_926 = 10'h39e == io_wrAddr_0 ? 2'h0 : lvtReg_926; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_927 = 10'h39f == io_wrAddr_0 ? 2'h0 : lvtReg_927; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_928 = 10'h3a0 == io_wrAddr_0 ? 2'h0 : lvtReg_928; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_929 = 10'h3a1 == io_wrAddr_0 ? 2'h0 : lvtReg_929; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_930 = 10'h3a2 == io_wrAddr_0 ? 2'h0 : lvtReg_930; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_931 = 10'h3a3 == io_wrAddr_0 ? 2'h0 : lvtReg_931; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_932 = 10'h3a4 == io_wrAddr_0 ? 2'h0 : lvtReg_932; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_933 = 10'h3a5 == io_wrAddr_0 ? 2'h0 : lvtReg_933; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_934 = 10'h3a6 == io_wrAddr_0 ? 2'h0 : lvtReg_934; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_935 = 10'h3a7 == io_wrAddr_0 ? 2'h0 : lvtReg_935; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_936 = 10'h3a8 == io_wrAddr_0 ? 2'h0 : lvtReg_936; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_937 = 10'h3a9 == io_wrAddr_0 ? 2'h0 : lvtReg_937; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_938 = 10'h3aa == io_wrAddr_0 ? 2'h0 : lvtReg_938; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_939 = 10'h3ab == io_wrAddr_0 ? 2'h0 : lvtReg_939; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_940 = 10'h3ac == io_wrAddr_0 ? 2'h0 : lvtReg_940; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_941 = 10'h3ad == io_wrAddr_0 ? 2'h0 : lvtReg_941; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_942 = 10'h3ae == io_wrAddr_0 ? 2'h0 : lvtReg_942; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_943 = 10'h3af == io_wrAddr_0 ? 2'h0 : lvtReg_943; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_944 = 10'h3b0 == io_wrAddr_0 ? 2'h0 : lvtReg_944; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_945 = 10'h3b1 == io_wrAddr_0 ? 2'h0 : lvtReg_945; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_946 = 10'h3b2 == io_wrAddr_0 ? 2'h0 : lvtReg_946; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_947 = 10'h3b3 == io_wrAddr_0 ? 2'h0 : lvtReg_947; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_948 = 10'h3b4 == io_wrAddr_0 ? 2'h0 : lvtReg_948; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_949 = 10'h3b5 == io_wrAddr_0 ? 2'h0 : lvtReg_949; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_950 = 10'h3b6 == io_wrAddr_0 ? 2'h0 : lvtReg_950; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_951 = 10'h3b7 == io_wrAddr_0 ? 2'h0 : lvtReg_951; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_952 = 10'h3b8 == io_wrAddr_0 ? 2'h0 : lvtReg_952; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_953 = 10'h3b9 == io_wrAddr_0 ? 2'h0 : lvtReg_953; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_954 = 10'h3ba == io_wrAddr_0 ? 2'h0 : lvtReg_954; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_955 = 10'h3bb == io_wrAddr_0 ? 2'h0 : lvtReg_955; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_956 = 10'h3bc == io_wrAddr_0 ? 2'h0 : lvtReg_956; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_957 = 10'h3bd == io_wrAddr_0 ? 2'h0 : lvtReg_957; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_958 = 10'h3be == io_wrAddr_0 ? 2'h0 : lvtReg_958; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_959 = 10'h3bf == io_wrAddr_0 ? 2'h0 : lvtReg_959; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_960 = 10'h3c0 == io_wrAddr_0 ? 2'h0 : lvtReg_960; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_961 = 10'h3c1 == io_wrAddr_0 ? 2'h0 : lvtReg_961; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_962 = 10'h3c2 == io_wrAddr_0 ? 2'h0 : lvtReg_962; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_963 = 10'h3c3 == io_wrAddr_0 ? 2'h0 : lvtReg_963; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_964 = 10'h3c4 == io_wrAddr_0 ? 2'h0 : lvtReg_964; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_965 = 10'h3c5 == io_wrAddr_0 ? 2'h0 : lvtReg_965; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_966 = 10'h3c6 == io_wrAddr_0 ? 2'h0 : lvtReg_966; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_967 = 10'h3c7 == io_wrAddr_0 ? 2'h0 : lvtReg_967; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_968 = 10'h3c8 == io_wrAddr_0 ? 2'h0 : lvtReg_968; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_969 = 10'h3c9 == io_wrAddr_0 ? 2'h0 : lvtReg_969; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_970 = 10'h3ca == io_wrAddr_0 ? 2'h0 : lvtReg_970; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_971 = 10'h3cb == io_wrAddr_0 ? 2'h0 : lvtReg_971; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_972 = 10'h3cc == io_wrAddr_0 ? 2'h0 : lvtReg_972; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_973 = 10'h3cd == io_wrAddr_0 ? 2'h0 : lvtReg_973; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_974 = 10'h3ce == io_wrAddr_0 ? 2'h0 : lvtReg_974; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_975 = 10'h3cf == io_wrAddr_0 ? 2'h0 : lvtReg_975; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_976 = 10'h3d0 == io_wrAddr_0 ? 2'h0 : lvtReg_976; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_977 = 10'h3d1 == io_wrAddr_0 ? 2'h0 : lvtReg_977; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_978 = 10'h3d2 == io_wrAddr_0 ? 2'h0 : lvtReg_978; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_979 = 10'h3d3 == io_wrAddr_0 ? 2'h0 : lvtReg_979; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_980 = 10'h3d4 == io_wrAddr_0 ? 2'h0 : lvtReg_980; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_981 = 10'h3d5 == io_wrAddr_0 ? 2'h0 : lvtReg_981; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_982 = 10'h3d6 == io_wrAddr_0 ? 2'h0 : lvtReg_982; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_983 = 10'h3d7 == io_wrAddr_0 ? 2'h0 : lvtReg_983; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_984 = 10'h3d8 == io_wrAddr_0 ? 2'h0 : lvtReg_984; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_985 = 10'h3d9 == io_wrAddr_0 ? 2'h0 : lvtReg_985; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_986 = 10'h3da == io_wrAddr_0 ? 2'h0 : lvtReg_986; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_987 = 10'h3db == io_wrAddr_0 ? 2'h0 : lvtReg_987; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_988 = 10'h3dc == io_wrAddr_0 ? 2'h0 : lvtReg_988; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_989 = 10'h3dd == io_wrAddr_0 ? 2'h0 : lvtReg_989; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_990 = 10'h3de == io_wrAddr_0 ? 2'h0 : lvtReg_990; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_991 = 10'h3df == io_wrAddr_0 ? 2'h0 : lvtReg_991; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_992 = 10'h3e0 == io_wrAddr_0 ? 2'h0 : lvtReg_992; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_993 = 10'h3e1 == io_wrAddr_0 ? 2'h0 : lvtReg_993; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_994 = 10'h3e2 == io_wrAddr_0 ? 2'h0 : lvtReg_994; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_995 = 10'h3e3 == io_wrAddr_0 ? 2'h0 : lvtReg_995; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_996 = 10'h3e4 == io_wrAddr_0 ? 2'h0 : lvtReg_996; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_997 = 10'h3e5 == io_wrAddr_0 ? 2'h0 : lvtReg_997; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_998 = 10'h3e6 == io_wrAddr_0 ? 2'h0 : lvtReg_998; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_999 = 10'h3e7 == io_wrAddr_0 ? 2'h0 : lvtReg_999; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1000 = 10'h3e8 == io_wrAddr_0 ? 2'h0 : lvtReg_1000; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1001 = 10'h3e9 == io_wrAddr_0 ? 2'h0 : lvtReg_1001; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1002 = 10'h3ea == io_wrAddr_0 ? 2'h0 : lvtReg_1002; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1003 = 10'h3eb == io_wrAddr_0 ? 2'h0 : lvtReg_1003; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1004 = 10'h3ec == io_wrAddr_0 ? 2'h0 : lvtReg_1004; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1005 = 10'h3ed == io_wrAddr_0 ? 2'h0 : lvtReg_1005; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1006 = 10'h3ee == io_wrAddr_0 ? 2'h0 : lvtReg_1006; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1007 = 10'h3ef == io_wrAddr_0 ? 2'h0 : lvtReg_1007; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1008 = 10'h3f0 == io_wrAddr_0 ? 2'h0 : lvtReg_1008; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1009 = 10'h3f1 == io_wrAddr_0 ? 2'h0 : lvtReg_1009; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1010 = 10'h3f2 == io_wrAddr_0 ? 2'h0 : lvtReg_1010; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1011 = 10'h3f3 == io_wrAddr_0 ? 2'h0 : lvtReg_1011; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1012 = 10'h3f4 == io_wrAddr_0 ? 2'h0 : lvtReg_1012; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1013 = 10'h3f5 == io_wrAddr_0 ? 2'h0 : lvtReg_1013; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1014 = 10'h3f6 == io_wrAddr_0 ? 2'h0 : lvtReg_1014; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1015 = 10'h3f7 == io_wrAddr_0 ? 2'h0 : lvtReg_1015; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1016 = 10'h3f8 == io_wrAddr_0 ? 2'h0 : lvtReg_1016; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1017 = 10'h3f9 == io_wrAddr_0 ? 2'h0 : lvtReg_1017; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1018 = 10'h3fa == io_wrAddr_0 ? 2'h0 : lvtReg_1018; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1019 = 10'h3fb == io_wrAddr_0 ? 2'h0 : lvtReg_1019; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1020 = 10'h3fc == io_wrAddr_0 ? 2'h0 : lvtReg_1020; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1021 = 10'h3fd == io_wrAddr_0 ? 2'h0 : lvtReg_1021; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1022 = 10'h3fe == io_wrAddr_0 ? 2'h0 : lvtReg_1022; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1023 = 10'h3ff == io_wrAddr_0 ? 2'h0 : lvtReg_1023; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1024 = io_wrEna_0 ? _GEN_0 : lvtReg_0; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1025 = io_wrEna_0 ? _GEN_1 : lvtReg_1; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1026 = io_wrEna_0 ? _GEN_2 : lvtReg_2; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1027 = io_wrEna_0 ? _GEN_3 : lvtReg_3; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1028 = io_wrEna_0 ? _GEN_4 : lvtReg_4; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1029 = io_wrEna_0 ? _GEN_5 : lvtReg_5; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1030 = io_wrEna_0 ? _GEN_6 : lvtReg_6; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1031 = io_wrEna_0 ? _GEN_7 : lvtReg_7; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1032 = io_wrEna_0 ? _GEN_8 : lvtReg_8; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1033 = io_wrEna_0 ? _GEN_9 : lvtReg_9; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1034 = io_wrEna_0 ? _GEN_10 : lvtReg_10; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1035 = io_wrEna_0 ? _GEN_11 : lvtReg_11; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1036 = io_wrEna_0 ? _GEN_12 : lvtReg_12; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1037 = io_wrEna_0 ? _GEN_13 : lvtReg_13; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1038 = io_wrEna_0 ? _GEN_14 : lvtReg_14; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1039 = io_wrEna_0 ? _GEN_15 : lvtReg_15; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1040 = io_wrEna_0 ? _GEN_16 : lvtReg_16; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1041 = io_wrEna_0 ? _GEN_17 : lvtReg_17; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1042 = io_wrEna_0 ? _GEN_18 : lvtReg_18; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1043 = io_wrEna_0 ? _GEN_19 : lvtReg_19; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1044 = io_wrEna_0 ? _GEN_20 : lvtReg_20; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1045 = io_wrEna_0 ? _GEN_21 : lvtReg_21; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1046 = io_wrEna_0 ? _GEN_22 : lvtReg_22; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1047 = io_wrEna_0 ? _GEN_23 : lvtReg_23; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1048 = io_wrEna_0 ? _GEN_24 : lvtReg_24; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1049 = io_wrEna_0 ? _GEN_25 : lvtReg_25; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1050 = io_wrEna_0 ? _GEN_26 : lvtReg_26; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1051 = io_wrEna_0 ? _GEN_27 : lvtReg_27; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1052 = io_wrEna_0 ? _GEN_28 : lvtReg_28; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1053 = io_wrEna_0 ? _GEN_29 : lvtReg_29; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1054 = io_wrEna_0 ? _GEN_30 : lvtReg_30; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1055 = io_wrEna_0 ? _GEN_31 : lvtReg_31; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1056 = io_wrEna_0 ? _GEN_32 : lvtReg_32; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1057 = io_wrEna_0 ? _GEN_33 : lvtReg_33; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1058 = io_wrEna_0 ? _GEN_34 : lvtReg_34; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1059 = io_wrEna_0 ? _GEN_35 : lvtReg_35; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1060 = io_wrEna_0 ? _GEN_36 : lvtReg_36; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1061 = io_wrEna_0 ? _GEN_37 : lvtReg_37; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1062 = io_wrEna_0 ? _GEN_38 : lvtReg_38; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1063 = io_wrEna_0 ? _GEN_39 : lvtReg_39; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1064 = io_wrEna_0 ? _GEN_40 : lvtReg_40; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1065 = io_wrEna_0 ? _GEN_41 : lvtReg_41; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1066 = io_wrEna_0 ? _GEN_42 : lvtReg_42; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1067 = io_wrEna_0 ? _GEN_43 : lvtReg_43; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1068 = io_wrEna_0 ? _GEN_44 : lvtReg_44; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1069 = io_wrEna_0 ? _GEN_45 : lvtReg_45; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1070 = io_wrEna_0 ? _GEN_46 : lvtReg_46; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1071 = io_wrEna_0 ? _GEN_47 : lvtReg_47; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1072 = io_wrEna_0 ? _GEN_48 : lvtReg_48; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1073 = io_wrEna_0 ? _GEN_49 : lvtReg_49; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1074 = io_wrEna_0 ? _GEN_50 : lvtReg_50; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1075 = io_wrEna_0 ? _GEN_51 : lvtReg_51; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1076 = io_wrEna_0 ? _GEN_52 : lvtReg_52; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1077 = io_wrEna_0 ? _GEN_53 : lvtReg_53; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1078 = io_wrEna_0 ? _GEN_54 : lvtReg_54; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1079 = io_wrEna_0 ? _GEN_55 : lvtReg_55; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1080 = io_wrEna_0 ? _GEN_56 : lvtReg_56; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1081 = io_wrEna_0 ? _GEN_57 : lvtReg_57; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1082 = io_wrEna_0 ? _GEN_58 : lvtReg_58; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1083 = io_wrEna_0 ? _GEN_59 : lvtReg_59; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1084 = io_wrEna_0 ? _GEN_60 : lvtReg_60; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1085 = io_wrEna_0 ? _GEN_61 : lvtReg_61; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1086 = io_wrEna_0 ? _GEN_62 : lvtReg_62; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1087 = io_wrEna_0 ? _GEN_63 : lvtReg_63; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1088 = io_wrEna_0 ? _GEN_64 : lvtReg_64; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1089 = io_wrEna_0 ? _GEN_65 : lvtReg_65; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1090 = io_wrEna_0 ? _GEN_66 : lvtReg_66; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1091 = io_wrEna_0 ? _GEN_67 : lvtReg_67; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1092 = io_wrEna_0 ? _GEN_68 : lvtReg_68; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1093 = io_wrEna_0 ? _GEN_69 : lvtReg_69; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1094 = io_wrEna_0 ? _GEN_70 : lvtReg_70; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1095 = io_wrEna_0 ? _GEN_71 : lvtReg_71; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1096 = io_wrEna_0 ? _GEN_72 : lvtReg_72; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1097 = io_wrEna_0 ? _GEN_73 : lvtReg_73; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1098 = io_wrEna_0 ? _GEN_74 : lvtReg_74; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1099 = io_wrEna_0 ? _GEN_75 : lvtReg_75; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1100 = io_wrEna_0 ? _GEN_76 : lvtReg_76; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1101 = io_wrEna_0 ? _GEN_77 : lvtReg_77; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1102 = io_wrEna_0 ? _GEN_78 : lvtReg_78; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1103 = io_wrEna_0 ? _GEN_79 : lvtReg_79; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1104 = io_wrEna_0 ? _GEN_80 : lvtReg_80; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1105 = io_wrEna_0 ? _GEN_81 : lvtReg_81; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1106 = io_wrEna_0 ? _GEN_82 : lvtReg_82; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1107 = io_wrEna_0 ? _GEN_83 : lvtReg_83; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1108 = io_wrEna_0 ? _GEN_84 : lvtReg_84; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1109 = io_wrEna_0 ? _GEN_85 : lvtReg_85; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1110 = io_wrEna_0 ? _GEN_86 : lvtReg_86; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1111 = io_wrEna_0 ? _GEN_87 : lvtReg_87; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1112 = io_wrEna_0 ? _GEN_88 : lvtReg_88; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1113 = io_wrEna_0 ? _GEN_89 : lvtReg_89; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1114 = io_wrEna_0 ? _GEN_90 : lvtReg_90; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1115 = io_wrEna_0 ? _GEN_91 : lvtReg_91; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1116 = io_wrEna_0 ? _GEN_92 : lvtReg_92; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1117 = io_wrEna_0 ? _GEN_93 : lvtReg_93; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1118 = io_wrEna_0 ? _GEN_94 : lvtReg_94; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1119 = io_wrEna_0 ? _GEN_95 : lvtReg_95; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1120 = io_wrEna_0 ? _GEN_96 : lvtReg_96; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1121 = io_wrEna_0 ? _GEN_97 : lvtReg_97; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1122 = io_wrEna_0 ? _GEN_98 : lvtReg_98; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1123 = io_wrEna_0 ? _GEN_99 : lvtReg_99; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1124 = io_wrEna_0 ? _GEN_100 : lvtReg_100; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1125 = io_wrEna_0 ? _GEN_101 : lvtReg_101; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1126 = io_wrEna_0 ? _GEN_102 : lvtReg_102; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1127 = io_wrEna_0 ? _GEN_103 : lvtReg_103; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1128 = io_wrEna_0 ? _GEN_104 : lvtReg_104; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1129 = io_wrEna_0 ? _GEN_105 : lvtReg_105; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1130 = io_wrEna_0 ? _GEN_106 : lvtReg_106; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1131 = io_wrEna_0 ? _GEN_107 : lvtReg_107; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1132 = io_wrEna_0 ? _GEN_108 : lvtReg_108; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1133 = io_wrEna_0 ? _GEN_109 : lvtReg_109; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1134 = io_wrEna_0 ? _GEN_110 : lvtReg_110; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1135 = io_wrEna_0 ? _GEN_111 : lvtReg_111; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1136 = io_wrEna_0 ? _GEN_112 : lvtReg_112; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1137 = io_wrEna_0 ? _GEN_113 : lvtReg_113; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1138 = io_wrEna_0 ? _GEN_114 : lvtReg_114; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1139 = io_wrEna_0 ? _GEN_115 : lvtReg_115; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1140 = io_wrEna_0 ? _GEN_116 : lvtReg_116; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1141 = io_wrEna_0 ? _GEN_117 : lvtReg_117; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1142 = io_wrEna_0 ? _GEN_118 : lvtReg_118; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1143 = io_wrEna_0 ? _GEN_119 : lvtReg_119; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1144 = io_wrEna_0 ? _GEN_120 : lvtReg_120; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1145 = io_wrEna_0 ? _GEN_121 : lvtReg_121; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1146 = io_wrEna_0 ? _GEN_122 : lvtReg_122; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1147 = io_wrEna_0 ? _GEN_123 : lvtReg_123; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1148 = io_wrEna_0 ? _GEN_124 : lvtReg_124; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1149 = io_wrEna_0 ? _GEN_125 : lvtReg_125; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1150 = io_wrEna_0 ? _GEN_126 : lvtReg_126; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1151 = io_wrEna_0 ? _GEN_127 : lvtReg_127; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1152 = io_wrEna_0 ? _GEN_128 : lvtReg_128; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1153 = io_wrEna_0 ? _GEN_129 : lvtReg_129; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1154 = io_wrEna_0 ? _GEN_130 : lvtReg_130; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1155 = io_wrEna_0 ? _GEN_131 : lvtReg_131; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1156 = io_wrEna_0 ? _GEN_132 : lvtReg_132; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1157 = io_wrEna_0 ? _GEN_133 : lvtReg_133; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1158 = io_wrEna_0 ? _GEN_134 : lvtReg_134; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1159 = io_wrEna_0 ? _GEN_135 : lvtReg_135; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1160 = io_wrEna_0 ? _GEN_136 : lvtReg_136; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1161 = io_wrEna_0 ? _GEN_137 : lvtReg_137; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1162 = io_wrEna_0 ? _GEN_138 : lvtReg_138; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1163 = io_wrEna_0 ? _GEN_139 : lvtReg_139; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1164 = io_wrEna_0 ? _GEN_140 : lvtReg_140; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1165 = io_wrEna_0 ? _GEN_141 : lvtReg_141; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1166 = io_wrEna_0 ? _GEN_142 : lvtReg_142; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1167 = io_wrEna_0 ? _GEN_143 : lvtReg_143; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1168 = io_wrEna_0 ? _GEN_144 : lvtReg_144; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1169 = io_wrEna_0 ? _GEN_145 : lvtReg_145; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1170 = io_wrEna_0 ? _GEN_146 : lvtReg_146; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1171 = io_wrEna_0 ? _GEN_147 : lvtReg_147; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1172 = io_wrEna_0 ? _GEN_148 : lvtReg_148; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1173 = io_wrEna_0 ? _GEN_149 : lvtReg_149; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1174 = io_wrEna_0 ? _GEN_150 : lvtReg_150; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1175 = io_wrEna_0 ? _GEN_151 : lvtReg_151; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1176 = io_wrEna_0 ? _GEN_152 : lvtReg_152; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1177 = io_wrEna_0 ? _GEN_153 : lvtReg_153; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1178 = io_wrEna_0 ? _GEN_154 : lvtReg_154; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1179 = io_wrEna_0 ? _GEN_155 : lvtReg_155; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1180 = io_wrEna_0 ? _GEN_156 : lvtReg_156; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1181 = io_wrEna_0 ? _GEN_157 : lvtReg_157; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1182 = io_wrEna_0 ? _GEN_158 : lvtReg_158; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1183 = io_wrEna_0 ? _GEN_159 : lvtReg_159; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1184 = io_wrEna_0 ? _GEN_160 : lvtReg_160; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1185 = io_wrEna_0 ? _GEN_161 : lvtReg_161; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1186 = io_wrEna_0 ? _GEN_162 : lvtReg_162; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1187 = io_wrEna_0 ? _GEN_163 : lvtReg_163; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1188 = io_wrEna_0 ? _GEN_164 : lvtReg_164; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1189 = io_wrEna_0 ? _GEN_165 : lvtReg_165; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1190 = io_wrEna_0 ? _GEN_166 : lvtReg_166; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1191 = io_wrEna_0 ? _GEN_167 : lvtReg_167; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1192 = io_wrEna_0 ? _GEN_168 : lvtReg_168; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1193 = io_wrEna_0 ? _GEN_169 : lvtReg_169; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1194 = io_wrEna_0 ? _GEN_170 : lvtReg_170; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1195 = io_wrEna_0 ? _GEN_171 : lvtReg_171; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1196 = io_wrEna_0 ? _GEN_172 : lvtReg_172; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1197 = io_wrEna_0 ? _GEN_173 : lvtReg_173; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1198 = io_wrEna_0 ? _GEN_174 : lvtReg_174; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1199 = io_wrEna_0 ? _GEN_175 : lvtReg_175; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1200 = io_wrEna_0 ? _GEN_176 : lvtReg_176; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1201 = io_wrEna_0 ? _GEN_177 : lvtReg_177; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1202 = io_wrEna_0 ? _GEN_178 : lvtReg_178; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1203 = io_wrEna_0 ? _GEN_179 : lvtReg_179; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1204 = io_wrEna_0 ? _GEN_180 : lvtReg_180; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1205 = io_wrEna_0 ? _GEN_181 : lvtReg_181; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1206 = io_wrEna_0 ? _GEN_182 : lvtReg_182; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1207 = io_wrEna_0 ? _GEN_183 : lvtReg_183; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1208 = io_wrEna_0 ? _GEN_184 : lvtReg_184; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1209 = io_wrEna_0 ? _GEN_185 : lvtReg_185; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1210 = io_wrEna_0 ? _GEN_186 : lvtReg_186; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1211 = io_wrEna_0 ? _GEN_187 : lvtReg_187; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1212 = io_wrEna_0 ? _GEN_188 : lvtReg_188; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1213 = io_wrEna_0 ? _GEN_189 : lvtReg_189; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1214 = io_wrEna_0 ? _GEN_190 : lvtReg_190; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1215 = io_wrEna_0 ? _GEN_191 : lvtReg_191; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1216 = io_wrEna_0 ? _GEN_192 : lvtReg_192; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1217 = io_wrEna_0 ? _GEN_193 : lvtReg_193; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1218 = io_wrEna_0 ? _GEN_194 : lvtReg_194; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1219 = io_wrEna_0 ? _GEN_195 : lvtReg_195; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1220 = io_wrEna_0 ? _GEN_196 : lvtReg_196; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1221 = io_wrEna_0 ? _GEN_197 : lvtReg_197; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1222 = io_wrEna_0 ? _GEN_198 : lvtReg_198; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1223 = io_wrEna_0 ? _GEN_199 : lvtReg_199; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1224 = io_wrEna_0 ? _GEN_200 : lvtReg_200; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1225 = io_wrEna_0 ? _GEN_201 : lvtReg_201; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1226 = io_wrEna_0 ? _GEN_202 : lvtReg_202; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1227 = io_wrEna_0 ? _GEN_203 : lvtReg_203; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1228 = io_wrEna_0 ? _GEN_204 : lvtReg_204; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1229 = io_wrEna_0 ? _GEN_205 : lvtReg_205; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1230 = io_wrEna_0 ? _GEN_206 : lvtReg_206; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1231 = io_wrEna_0 ? _GEN_207 : lvtReg_207; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1232 = io_wrEna_0 ? _GEN_208 : lvtReg_208; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1233 = io_wrEna_0 ? _GEN_209 : lvtReg_209; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1234 = io_wrEna_0 ? _GEN_210 : lvtReg_210; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1235 = io_wrEna_0 ? _GEN_211 : lvtReg_211; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1236 = io_wrEna_0 ? _GEN_212 : lvtReg_212; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1237 = io_wrEna_0 ? _GEN_213 : lvtReg_213; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1238 = io_wrEna_0 ? _GEN_214 : lvtReg_214; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1239 = io_wrEna_0 ? _GEN_215 : lvtReg_215; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1240 = io_wrEna_0 ? _GEN_216 : lvtReg_216; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1241 = io_wrEna_0 ? _GEN_217 : lvtReg_217; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1242 = io_wrEna_0 ? _GEN_218 : lvtReg_218; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1243 = io_wrEna_0 ? _GEN_219 : lvtReg_219; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1244 = io_wrEna_0 ? _GEN_220 : lvtReg_220; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1245 = io_wrEna_0 ? _GEN_221 : lvtReg_221; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1246 = io_wrEna_0 ? _GEN_222 : lvtReg_222; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1247 = io_wrEna_0 ? _GEN_223 : lvtReg_223; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1248 = io_wrEna_0 ? _GEN_224 : lvtReg_224; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1249 = io_wrEna_0 ? _GEN_225 : lvtReg_225; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1250 = io_wrEna_0 ? _GEN_226 : lvtReg_226; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1251 = io_wrEna_0 ? _GEN_227 : lvtReg_227; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1252 = io_wrEna_0 ? _GEN_228 : lvtReg_228; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1253 = io_wrEna_0 ? _GEN_229 : lvtReg_229; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1254 = io_wrEna_0 ? _GEN_230 : lvtReg_230; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1255 = io_wrEna_0 ? _GEN_231 : lvtReg_231; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1256 = io_wrEna_0 ? _GEN_232 : lvtReg_232; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1257 = io_wrEna_0 ? _GEN_233 : lvtReg_233; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1258 = io_wrEna_0 ? _GEN_234 : lvtReg_234; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1259 = io_wrEna_0 ? _GEN_235 : lvtReg_235; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1260 = io_wrEna_0 ? _GEN_236 : lvtReg_236; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1261 = io_wrEna_0 ? _GEN_237 : lvtReg_237; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1262 = io_wrEna_0 ? _GEN_238 : lvtReg_238; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1263 = io_wrEna_0 ? _GEN_239 : lvtReg_239; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1264 = io_wrEna_0 ? _GEN_240 : lvtReg_240; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1265 = io_wrEna_0 ? _GEN_241 : lvtReg_241; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1266 = io_wrEna_0 ? _GEN_242 : lvtReg_242; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1267 = io_wrEna_0 ? _GEN_243 : lvtReg_243; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1268 = io_wrEna_0 ? _GEN_244 : lvtReg_244; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1269 = io_wrEna_0 ? _GEN_245 : lvtReg_245; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1270 = io_wrEna_0 ? _GEN_246 : lvtReg_246; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1271 = io_wrEna_0 ? _GEN_247 : lvtReg_247; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1272 = io_wrEna_0 ? _GEN_248 : lvtReg_248; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1273 = io_wrEna_0 ? _GEN_249 : lvtReg_249; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1274 = io_wrEna_0 ? _GEN_250 : lvtReg_250; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1275 = io_wrEna_0 ? _GEN_251 : lvtReg_251; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1276 = io_wrEna_0 ? _GEN_252 : lvtReg_252; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1277 = io_wrEna_0 ? _GEN_253 : lvtReg_253; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1278 = io_wrEna_0 ? _GEN_254 : lvtReg_254; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1279 = io_wrEna_0 ? _GEN_255 : lvtReg_255; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1280 = io_wrEna_0 ? _GEN_256 : lvtReg_256; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1281 = io_wrEna_0 ? _GEN_257 : lvtReg_257; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1282 = io_wrEna_0 ? _GEN_258 : lvtReg_258; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1283 = io_wrEna_0 ? _GEN_259 : lvtReg_259; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1284 = io_wrEna_0 ? _GEN_260 : lvtReg_260; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1285 = io_wrEna_0 ? _GEN_261 : lvtReg_261; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1286 = io_wrEna_0 ? _GEN_262 : lvtReg_262; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1287 = io_wrEna_0 ? _GEN_263 : lvtReg_263; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1288 = io_wrEna_0 ? _GEN_264 : lvtReg_264; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1289 = io_wrEna_0 ? _GEN_265 : lvtReg_265; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1290 = io_wrEna_0 ? _GEN_266 : lvtReg_266; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1291 = io_wrEna_0 ? _GEN_267 : lvtReg_267; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1292 = io_wrEna_0 ? _GEN_268 : lvtReg_268; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1293 = io_wrEna_0 ? _GEN_269 : lvtReg_269; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1294 = io_wrEna_0 ? _GEN_270 : lvtReg_270; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1295 = io_wrEna_0 ? _GEN_271 : lvtReg_271; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1296 = io_wrEna_0 ? _GEN_272 : lvtReg_272; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1297 = io_wrEna_0 ? _GEN_273 : lvtReg_273; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1298 = io_wrEna_0 ? _GEN_274 : lvtReg_274; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1299 = io_wrEna_0 ? _GEN_275 : lvtReg_275; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1300 = io_wrEna_0 ? _GEN_276 : lvtReg_276; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1301 = io_wrEna_0 ? _GEN_277 : lvtReg_277; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1302 = io_wrEna_0 ? _GEN_278 : lvtReg_278; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1303 = io_wrEna_0 ? _GEN_279 : lvtReg_279; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1304 = io_wrEna_0 ? _GEN_280 : lvtReg_280; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1305 = io_wrEna_0 ? _GEN_281 : lvtReg_281; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1306 = io_wrEna_0 ? _GEN_282 : lvtReg_282; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1307 = io_wrEna_0 ? _GEN_283 : lvtReg_283; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1308 = io_wrEna_0 ? _GEN_284 : lvtReg_284; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1309 = io_wrEna_0 ? _GEN_285 : lvtReg_285; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1310 = io_wrEna_0 ? _GEN_286 : lvtReg_286; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1311 = io_wrEna_0 ? _GEN_287 : lvtReg_287; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1312 = io_wrEna_0 ? _GEN_288 : lvtReg_288; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1313 = io_wrEna_0 ? _GEN_289 : lvtReg_289; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1314 = io_wrEna_0 ? _GEN_290 : lvtReg_290; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1315 = io_wrEna_0 ? _GEN_291 : lvtReg_291; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1316 = io_wrEna_0 ? _GEN_292 : lvtReg_292; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1317 = io_wrEna_0 ? _GEN_293 : lvtReg_293; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1318 = io_wrEna_0 ? _GEN_294 : lvtReg_294; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1319 = io_wrEna_0 ? _GEN_295 : lvtReg_295; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1320 = io_wrEna_0 ? _GEN_296 : lvtReg_296; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1321 = io_wrEna_0 ? _GEN_297 : lvtReg_297; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1322 = io_wrEna_0 ? _GEN_298 : lvtReg_298; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1323 = io_wrEna_0 ? _GEN_299 : lvtReg_299; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1324 = io_wrEna_0 ? _GEN_300 : lvtReg_300; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1325 = io_wrEna_0 ? _GEN_301 : lvtReg_301; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1326 = io_wrEna_0 ? _GEN_302 : lvtReg_302; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1327 = io_wrEna_0 ? _GEN_303 : lvtReg_303; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1328 = io_wrEna_0 ? _GEN_304 : lvtReg_304; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1329 = io_wrEna_0 ? _GEN_305 : lvtReg_305; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1330 = io_wrEna_0 ? _GEN_306 : lvtReg_306; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1331 = io_wrEna_0 ? _GEN_307 : lvtReg_307; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1332 = io_wrEna_0 ? _GEN_308 : lvtReg_308; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1333 = io_wrEna_0 ? _GEN_309 : lvtReg_309; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1334 = io_wrEna_0 ? _GEN_310 : lvtReg_310; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1335 = io_wrEna_0 ? _GEN_311 : lvtReg_311; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1336 = io_wrEna_0 ? _GEN_312 : lvtReg_312; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1337 = io_wrEna_0 ? _GEN_313 : lvtReg_313; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1338 = io_wrEna_0 ? _GEN_314 : lvtReg_314; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1339 = io_wrEna_0 ? _GEN_315 : lvtReg_315; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1340 = io_wrEna_0 ? _GEN_316 : lvtReg_316; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1341 = io_wrEna_0 ? _GEN_317 : lvtReg_317; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1342 = io_wrEna_0 ? _GEN_318 : lvtReg_318; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1343 = io_wrEna_0 ? _GEN_319 : lvtReg_319; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1344 = io_wrEna_0 ? _GEN_320 : lvtReg_320; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1345 = io_wrEna_0 ? _GEN_321 : lvtReg_321; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1346 = io_wrEna_0 ? _GEN_322 : lvtReg_322; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1347 = io_wrEna_0 ? _GEN_323 : lvtReg_323; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1348 = io_wrEna_0 ? _GEN_324 : lvtReg_324; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1349 = io_wrEna_0 ? _GEN_325 : lvtReg_325; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1350 = io_wrEna_0 ? _GEN_326 : lvtReg_326; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1351 = io_wrEna_0 ? _GEN_327 : lvtReg_327; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1352 = io_wrEna_0 ? _GEN_328 : lvtReg_328; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1353 = io_wrEna_0 ? _GEN_329 : lvtReg_329; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1354 = io_wrEna_0 ? _GEN_330 : lvtReg_330; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1355 = io_wrEna_0 ? _GEN_331 : lvtReg_331; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1356 = io_wrEna_0 ? _GEN_332 : lvtReg_332; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1357 = io_wrEna_0 ? _GEN_333 : lvtReg_333; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1358 = io_wrEna_0 ? _GEN_334 : lvtReg_334; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1359 = io_wrEna_0 ? _GEN_335 : lvtReg_335; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1360 = io_wrEna_0 ? _GEN_336 : lvtReg_336; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1361 = io_wrEna_0 ? _GEN_337 : lvtReg_337; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1362 = io_wrEna_0 ? _GEN_338 : lvtReg_338; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1363 = io_wrEna_0 ? _GEN_339 : lvtReg_339; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1364 = io_wrEna_0 ? _GEN_340 : lvtReg_340; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1365 = io_wrEna_0 ? _GEN_341 : lvtReg_341; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1366 = io_wrEna_0 ? _GEN_342 : lvtReg_342; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1367 = io_wrEna_0 ? _GEN_343 : lvtReg_343; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1368 = io_wrEna_0 ? _GEN_344 : lvtReg_344; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1369 = io_wrEna_0 ? _GEN_345 : lvtReg_345; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1370 = io_wrEna_0 ? _GEN_346 : lvtReg_346; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1371 = io_wrEna_0 ? _GEN_347 : lvtReg_347; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1372 = io_wrEna_0 ? _GEN_348 : lvtReg_348; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1373 = io_wrEna_0 ? _GEN_349 : lvtReg_349; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1374 = io_wrEna_0 ? _GEN_350 : lvtReg_350; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1375 = io_wrEna_0 ? _GEN_351 : lvtReg_351; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1376 = io_wrEna_0 ? _GEN_352 : lvtReg_352; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1377 = io_wrEna_0 ? _GEN_353 : lvtReg_353; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1378 = io_wrEna_0 ? _GEN_354 : lvtReg_354; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1379 = io_wrEna_0 ? _GEN_355 : lvtReg_355; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1380 = io_wrEna_0 ? _GEN_356 : lvtReg_356; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1381 = io_wrEna_0 ? _GEN_357 : lvtReg_357; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1382 = io_wrEna_0 ? _GEN_358 : lvtReg_358; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1383 = io_wrEna_0 ? _GEN_359 : lvtReg_359; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1384 = io_wrEna_0 ? _GEN_360 : lvtReg_360; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1385 = io_wrEna_0 ? _GEN_361 : lvtReg_361; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1386 = io_wrEna_0 ? _GEN_362 : lvtReg_362; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1387 = io_wrEna_0 ? _GEN_363 : lvtReg_363; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1388 = io_wrEna_0 ? _GEN_364 : lvtReg_364; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1389 = io_wrEna_0 ? _GEN_365 : lvtReg_365; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1390 = io_wrEna_0 ? _GEN_366 : lvtReg_366; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1391 = io_wrEna_0 ? _GEN_367 : lvtReg_367; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1392 = io_wrEna_0 ? _GEN_368 : lvtReg_368; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1393 = io_wrEna_0 ? _GEN_369 : lvtReg_369; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1394 = io_wrEna_0 ? _GEN_370 : lvtReg_370; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1395 = io_wrEna_0 ? _GEN_371 : lvtReg_371; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1396 = io_wrEna_0 ? _GEN_372 : lvtReg_372; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1397 = io_wrEna_0 ? _GEN_373 : lvtReg_373; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1398 = io_wrEna_0 ? _GEN_374 : lvtReg_374; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1399 = io_wrEna_0 ? _GEN_375 : lvtReg_375; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1400 = io_wrEna_0 ? _GEN_376 : lvtReg_376; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1401 = io_wrEna_0 ? _GEN_377 : lvtReg_377; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1402 = io_wrEna_0 ? _GEN_378 : lvtReg_378; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1403 = io_wrEna_0 ? _GEN_379 : lvtReg_379; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1404 = io_wrEna_0 ? _GEN_380 : lvtReg_380; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1405 = io_wrEna_0 ? _GEN_381 : lvtReg_381; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1406 = io_wrEna_0 ? _GEN_382 : lvtReg_382; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1407 = io_wrEna_0 ? _GEN_383 : lvtReg_383; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1408 = io_wrEna_0 ? _GEN_384 : lvtReg_384; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1409 = io_wrEna_0 ? _GEN_385 : lvtReg_385; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1410 = io_wrEna_0 ? _GEN_386 : lvtReg_386; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1411 = io_wrEna_0 ? _GEN_387 : lvtReg_387; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1412 = io_wrEna_0 ? _GEN_388 : lvtReg_388; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1413 = io_wrEna_0 ? _GEN_389 : lvtReg_389; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1414 = io_wrEna_0 ? _GEN_390 : lvtReg_390; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1415 = io_wrEna_0 ? _GEN_391 : lvtReg_391; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1416 = io_wrEna_0 ? _GEN_392 : lvtReg_392; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1417 = io_wrEna_0 ? _GEN_393 : lvtReg_393; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1418 = io_wrEna_0 ? _GEN_394 : lvtReg_394; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1419 = io_wrEna_0 ? _GEN_395 : lvtReg_395; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1420 = io_wrEna_0 ? _GEN_396 : lvtReg_396; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1421 = io_wrEna_0 ? _GEN_397 : lvtReg_397; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1422 = io_wrEna_0 ? _GEN_398 : lvtReg_398; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1423 = io_wrEna_0 ? _GEN_399 : lvtReg_399; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1424 = io_wrEna_0 ? _GEN_400 : lvtReg_400; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1425 = io_wrEna_0 ? _GEN_401 : lvtReg_401; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1426 = io_wrEna_0 ? _GEN_402 : lvtReg_402; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1427 = io_wrEna_0 ? _GEN_403 : lvtReg_403; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1428 = io_wrEna_0 ? _GEN_404 : lvtReg_404; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1429 = io_wrEna_0 ? _GEN_405 : lvtReg_405; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1430 = io_wrEna_0 ? _GEN_406 : lvtReg_406; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1431 = io_wrEna_0 ? _GEN_407 : lvtReg_407; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1432 = io_wrEna_0 ? _GEN_408 : lvtReg_408; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1433 = io_wrEna_0 ? _GEN_409 : lvtReg_409; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1434 = io_wrEna_0 ? _GEN_410 : lvtReg_410; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1435 = io_wrEna_0 ? _GEN_411 : lvtReg_411; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1436 = io_wrEna_0 ? _GEN_412 : lvtReg_412; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1437 = io_wrEna_0 ? _GEN_413 : lvtReg_413; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1438 = io_wrEna_0 ? _GEN_414 : lvtReg_414; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1439 = io_wrEna_0 ? _GEN_415 : lvtReg_415; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1440 = io_wrEna_0 ? _GEN_416 : lvtReg_416; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1441 = io_wrEna_0 ? _GEN_417 : lvtReg_417; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1442 = io_wrEna_0 ? _GEN_418 : lvtReg_418; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1443 = io_wrEna_0 ? _GEN_419 : lvtReg_419; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1444 = io_wrEna_0 ? _GEN_420 : lvtReg_420; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1445 = io_wrEna_0 ? _GEN_421 : lvtReg_421; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1446 = io_wrEna_0 ? _GEN_422 : lvtReg_422; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1447 = io_wrEna_0 ? _GEN_423 : lvtReg_423; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1448 = io_wrEna_0 ? _GEN_424 : lvtReg_424; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1449 = io_wrEna_0 ? _GEN_425 : lvtReg_425; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1450 = io_wrEna_0 ? _GEN_426 : lvtReg_426; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1451 = io_wrEna_0 ? _GEN_427 : lvtReg_427; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1452 = io_wrEna_0 ? _GEN_428 : lvtReg_428; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1453 = io_wrEna_0 ? _GEN_429 : lvtReg_429; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1454 = io_wrEna_0 ? _GEN_430 : lvtReg_430; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1455 = io_wrEna_0 ? _GEN_431 : lvtReg_431; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1456 = io_wrEna_0 ? _GEN_432 : lvtReg_432; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1457 = io_wrEna_0 ? _GEN_433 : lvtReg_433; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1458 = io_wrEna_0 ? _GEN_434 : lvtReg_434; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1459 = io_wrEna_0 ? _GEN_435 : lvtReg_435; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1460 = io_wrEna_0 ? _GEN_436 : lvtReg_436; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1461 = io_wrEna_0 ? _GEN_437 : lvtReg_437; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1462 = io_wrEna_0 ? _GEN_438 : lvtReg_438; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1463 = io_wrEna_0 ? _GEN_439 : lvtReg_439; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1464 = io_wrEna_0 ? _GEN_440 : lvtReg_440; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1465 = io_wrEna_0 ? _GEN_441 : lvtReg_441; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1466 = io_wrEna_0 ? _GEN_442 : lvtReg_442; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1467 = io_wrEna_0 ? _GEN_443 : lvtReg_443; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1468 = io_wrEna_0 ? _GEN_444 : lvtReg_444; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1469 = io_wrEna_0 ? _GEN_445 : lvtReg_445; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1470 = io_wrEna_0 ? _GEN_446 : lvtReg_446; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1471 = io_wrEna_0 ? _GEN_447 : lvtReg_447; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1472 = io_wrEna_0 ? _GEN_448 : lvtReg_448; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1473 = io_wrEna_0 ? _GEN_449 : lvtReg_449; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1474 = io_wrEna_0 ? _GEN_450 : lvtReg_450; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1475 = io_wrEna_0 ? _GEN_451 : lvtReg_451; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1476 = io_wrEna_0 ? _GEN_452 : lvtReg_452; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1477 = io_wrEna_0 ? _GEN_453 : lvtReg_453; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1478 = io_wrEna_0 ? _GEN_454 : lvtReg_454; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1479 = io_wrEna_0 ? _GEN_455 : lvtReg_455; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1480 = io_wrEna_0 ? _GEN_456 : lvtReg_456; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1481 = io_wrEna_0 ? _GEN_457 : lvtReg_457; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1482 = io_wrEna_0 ? _GEN_458 : lvtReg_458; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1483 = io_wrEna_0 ? _GEN_459 : lvtReg_459; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1484 = io_wrEna_0 ? _GEN_460 : lvtReg_460; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1485 = io_wrEna_0 ? _GEN_461 : lvtReg_461; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1486 = io_wrEna_0 ? _GEN_462 : lvtReg_462; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1487 = io_wrEna_0 ? _GEN_463 : lvtReg_463; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1488 = io_wrEna_0 ? _GEN_464 : lvtReg_464; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1489 = io_wrEna_0 ? _GEN_465 : lvtReg_465; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1490 = io_wrEna_0 ? _GEN_466 : lvtReg_466; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1491 = io_wrEna_0 ? _GEN_467 : lvtReg_467; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1492 = io_wrEna_0 ? _GEN_468 : lvtReg_468; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1493 = io_wrEna_0 ? _GEN_469 : lvtReg_469; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1494 = io_wrEna_0 ? _GEN_470 : lvtReg_470; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1495 = io_wrEna_0 ? _GEN_471 : lvtReg_471; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1496 = io_wrEna_0 ? _GEN_472 : lvtReg_472; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1497 = io_wrEna_0 ? _GEN_473 : lvtReg_473; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1498 = io_wrEna_0 ? _GEN_474 : lvtReg_474; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1499 = io_wrEna_0 ? _GEN_475 : lvtReg_475; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1500 = io_wrEna_0 ? _GEN_476 : lvtReg_476; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1501 = io_wrEna_0 ? _GEN_477 : lvtReg_477; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1502 = io_wrEna_0 ? _GEN_478 : lvtReg_478; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1503 = io_wrEna_0 ? _GEN_479 : lvtReg_479; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1504 = io_wrEna_0 ? _GEN_480 : lvtReg_480; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1505 = io_wrEna_0 ? _GEN_481 : lvtReg_481; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1506 = io_wrEna_0 ? _GEN_482 : lvtReg_482; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1507 = io_wrEna_0 ? _GEN_483 : lvtReg_483; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1508 = io_wrEna_0 ? _GEN_484 : lvtReg_484; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1509 = io_wrEna_0 ? _GEN_485 : lvtReg_485; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1510 = io_wrEna_0 ? _GEN_486 : lvtReg_486; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1511 = io_wrEna_0 ? _GEN_487 : lvtReg_487; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1512 = io_wrEna_0 ? _GEN_488 : lvtReg_488; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1513 = io_wrEna_0 ? _GEN_489 : lvtReg_489; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1514 = io_wrEna_0 ? _GEN_490 : lvtReg_490; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1515 = io_wrEna_0 ? _GEN_491 : lvtReg_491; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1516 = io_wrEna_0 ? _GEN_492 : lvtReg_492; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1517 = io_wrEna_0 ? _GEN_493 : lvtReg_493; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1518 = io_wrEna_0 ? _GEN_494 : lvtReg_494; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1519 = io_wrEna_0 ? _GEN_495 : lvtReg_495; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1520 = io_wrEna_0 ? _GEN_496 : lvtReg_496; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1521 = io_wrEna_0 ? _GEN_497 : lvtReg_497; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1522 = io_wrEna_0 ? _GEN_498 : lvtReg_498; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1523 = io_wrEna_0 ? _GEN_499 : lvtReg_499; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1524 = io_wrEna_0 ? _GEN_500 : lvtReg_500; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1525 = io_wrEna_0 ? _GEN_501 : lvtReg_501; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1526 = io_wrEna_0 ? _GEN_502 : lvtReg_502; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1527 = io_wrEna_0 ? _GEN_503 : lvtReg_503; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1528 = io_wrEna_0 ? _GEN_504 : lvtReg_504; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1529 = io_wrEna_0 ? _GEN_505 : lvtReg_505; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1530 = io_wrEna_0 ? _GEN_506 : lvtReg_506; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1531 = io_wrEna_0 ? _GEN_507 : lvtReg_507; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1532 = io_wrEna_0 ? _GEN_508 : lvtReg_508; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1533 = io_wrEna_0 ? _GEN_509 : lvtReg_509; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1534 = io_wrEna_0 ? _GEN_510 : lvtReg_510; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1535 = io_wrEna_0 ? _GEN_511 : lvtReg_511; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1536 = io_wrEna_0 ? _GEN_512 : lvtReg_512; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1537 = io_wrEna_0 ? _GEN_513 : lvtReg_513; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1538 = io_wrEna_0 ? _GEN_514 : lvtReg_514; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1539 = io_wrEna_0 ? _GEN_515 : lvtReg_515; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1540 = io_wrEna_0 ? _GEN_516 : lvtReg_516; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1541 = io_wrEna_0 ? _GEN_517 : lvtReg_517; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1542 = io_wrEna_0 ? _GEN_518 : lvtReg_518; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1543 = io_wrEna_0 ? _GEN_519 : lvtReg_519; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1544 = io_wrEna_0 ? _GEN_520 : lvtReg_520; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1545 = io_wrEna_0 ? _GEN_521 : lvtReg_521; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1546 = io_wrEna_0 ? _GEN_522 : lvtReg_522; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1547 = io_wrEna_0 ? _GEN_523 : lvtReg_523; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1548 = io_wrEna_0 ? _GEN_524 : lvtReg_524; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1549 = io_wrEna_0 ? _GEN_525 : lvtReg_525; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1550 = io_wrEna_0 ? _GEN_526 : lvtReg_526; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1551 = io_wrEna_0 ? _GEN_527 : lvtReg_527; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1552 = io_wrEna_0 ? _GEN_528 : lvtReg_528; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1553 = io_wrEna_0 ? _GEN_529 : lvtReg_529; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1554 = io_wrEna_0 ? _GEN_530 : lvtReg_530; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1555 = io_wrEna_0 ? _GEN_531 : lvtReg_531; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1556 = io_wrEna_0 ? _GEN_532 : lvtReg_532; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1557 = io_wrEna_0 ? _GEN_533 : lvtReg_533; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1558 = io_wrEna_0 ? _GEN_534 : lvtReg_534; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1559 = io_wrEna_0 ? _GEN_535 : lvtReg_535; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1560 = io_wrEna_0 ? _GEN_536 : lvtReg_536; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1561 = io_wrEna_0 ? _GEN_537 : lvtReg_537; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1562 = io_wrEna_0 ? _GEN_538 : lvtReg_538; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1563 = io_wrEna_0 ? _GEN_539 : lvtReg_539; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1564 = io_wrEna_0 ? _GEN_540 : lvtReg_540; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1565 = io_wrEna_0 ? _GEN_541 : lvtReg_541; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1566 = io_wrEna_0 ? _GEN_542 : lvtReg_542; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1567 = io_wrEna_0 ? _GEN_543 : lvtReg_543; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1568 = io_wrEna_0 ? _GEN_544 : lvtReg_544; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1569 = io_wrEna_0 ? _GEN_545 : lvtReg_545; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1570 = io_wrEna_0 ? _GEN_546 : lvtReg_546; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1571 = io_wrEna_0 ? _GEN_547 : lvtReg_547; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1572 = io_wrEna_0 ? _GEN_548 : lvtReg_548; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1573 = io_wrEna_0 ? _GEN_549 : lvtReg_549; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1574 = io_wrEna_0 ? _GEN_550 : lvtReg_550; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1575 = io_wrEna_0 ? _GEN_551 : lvtReg_551; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1576 = io_wrEna_0 ? _GEN_552 : lvtReg_552; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1577 = io_wrEna_0 ? _GEN_553 : lvtReg_553; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1578 = io_wrEna_0 ? _GEN_554 : lvtReg_554; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1579 = io_wrEna_0 ? _GEN_555 : lvtReg_555; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1580 = io_wrEna_0 ? _GEN_556 : lvtReg_556; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1581 = io_wrEna_0 ? _GEN_557 : lvtReg_557; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1582 = io_wrEna_0 ? _GEN_558 : lvtReg_558; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1583 = io_wrEna_0 ? _GEN_559 : lvtReg_559; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1584 = io_wrEna_0 ? _GEN_560 : lvtReg_560; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1585 = io_wrEna_0 ? _GEN_561 : lvtReg_561; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1586 = io_wrEna_0 ? _GEN_562 : lvtReg_562; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1587 = io_wrEna_0 ? _GEN_563 : lvtReg_563; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1588 = io_wrEna_0 ? _GEN_564 : lvtReg_564; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1589 = io_wrEna_0 ? _GEN_565 : lvtReg_565; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1590 = io_wrEna_0 ? _GEN_566 : lvtReg_566; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1591 = io_wrEna_0 ? _GEN_567 : lvtReg_567; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1592 = io_wrEna_0 ? _GEN_568 : lvtReg_568; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1593 = io_wrEna_0 ? _GEN_569 : lvtReg_569; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1594 = io_wrEna_0 ? _GEN_570 : lvtReg_570; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1595 = io_wrEna_0 ? _GEN_571 : lvtReg_571; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1596 = io_wrEna_0 ? _GEN_572 : lvtReg_572; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1597 = io_wrEna_0 ? _GEN_573 : lvtReg_573; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1598 = io_wrEna_0 ? _GEN_574 : lvtReg_574; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1599 = io_wrEna_0 ? _GEN_575 : lvtReg_575; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1600 = io_wrEna_0 ? _GEN_576 : lvtReg_576; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1601 = io_wrEna_0 ? _GEN_577 : lvtReg_577; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1602 = io_wrEna_0 ? _GEN_578 : lvtReg_578; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1603 = io_wrEna_0 ? _GEN_579 : lvtReg_579; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1604 = io_wrEna_0 ? _GEN_580 : lvtReg_580; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1605 = io_wrEna_0 ? _GEN_581 : lvtReg_581; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1606 = io_wrEna_0 ? _GEN_582 : lvtReg_582; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1607 = io_wrEna_0 ? _GEN_583 : lvtReg_583; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1608 = io_wrEna_0 ? _GEN_584 : lvtReg_584; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1609 = io_wrEna_0 ? _GEN_585 : lvtReg_585; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1610 = io_wrEna_0 ? _GEN_586 : lvtReg_586; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1611 = io_wrEna_0 ? _GEN_587 : lvtReg_587; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1612 = io_wrEna_0 ? _GEN_588 : lvtReg_588; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1613 = io_wrEna_0 ? _GEN_589 : lvtReg_589; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1614 = io_wrEna_0 ? _GEN_590 : lvtReg_590; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1615 = io_wrEna_0 ? _GEN_591 : lvtReg_591; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1616 = io_wrEna_0 ? _GEN_592 : lvtReg_592; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1617 = io_wrEna_0 ? _GEN_593 : lvtReg_593; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1618 = io_wrEna_0 ? _GEN_594 : lvtReg_594; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1619 = io_wrEna_0 ? _GEN_595 : lvtReg_595; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1620 = io_wrEna_0 ? _GEN_596 : lvtReg_596; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1621 = io_wrEna_0 ? _GEN_597 : lvtReg_597; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1622 = io_wrEna_0 ? _GEN_598 : lvtReg_598; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1623 = io_wrEna_0 ? _GEN_599 : lvtReg_599; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1624 = io_wrEna_0 ? _GEN_600 : lvtReg_600; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1625 = io_wrEna_0 ? _GEN_601 : lvtReg_601; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1626 = io_wrEna_0 ? _GEN_602 : lvtReg_602; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1627 = io_wrEna_0 ? _GEN_603 : lvtReg_603; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1628 = io_wrEna_0 ? _GEN_604 : lvtReg_604; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1629 = io_wrEna_0 ? _GEN_605 : lvtReg_605; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1630 = io_wrEna_0 ? _GEN_606 : lvtReg_606; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1631 = io_wrEna_0 ? _GEN_607 : lvtReg_607; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1632 = io_wrEna_0 ? _GEN_608 : lvtReg_608; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1633 = io_wrEna_0 ? _GEN_609 : lvtReg_609; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1634 = io_wrEna_0 ? _GEN_610 : lvtReg_610; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1635 = io_wrEna_0 ? _GEN_611 : lvtReg_611; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1636 = io_wrEna_0 ? _GEN_612 : lvtReg_612; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1637 = io_wrEna_0 ? _GEN_613 : lvtReg_613; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1638 = io_wrEna_0 ? _GEN_614 : lvtReg_614; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1639 = io_wrEna_0 ? _GEN_615 : lvtReg_615; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1640 = io_wrEna_0 ? _GEN_616 : lvtReg_616; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1641 = io_wrEna_0 ? _GEN_617 : lvtReg_617; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1642 = io_wrEna_0 ? _GEN_618 : lvtReg_618; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1643 = io_wrEna_0 ? _GEN_619 : lvtReg_619; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1644 = io_wrEna_0 ? _GEN_620 : lvtReg_620; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1645 = io_wrEna_0 ? _GEN_621 : lvtReg_621; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1646 = io_wrEna_0 ? _GEN_622 : lvtReg_622; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1647 = io_wrEna_0 ? _GEN_623 : lvtReg_623; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1648 = io_wrEna_0 ? _GEN_624 : lvtReg_624; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1649 = io_wrEna_0 ? _GEN_625 : lvtReg_625; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1650 = io_wrEna_0 ? _GEN_626 : lvtReg_626; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1651 = io_wrEna_0 ? _GEN_627 : lvtReg_627; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1652 = io_wrEna_0 ? _GEN_628 : lvtReg_628; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1653 = io_wrEna_0 ? _GEN_629 : lvtReg_629; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1654 = io_wrEna_0 ? _GEN_630 : lvtReg_630; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1655 = io_wrEna_0 ? _GEN_631 : lvtReg_631; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1656 = io_wrEna_0 ? _GEN_632 : lvtReg_632; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1657 = io_wrEna_0 ? _GEN_633 : lvtReg_633; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1658 = io_wrEna_0 ? _GEN_634 : lvtReg_634; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1659 = io_wrEna_0 ? _GEN_635 : lvtReg_635; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1660 = io_wrEna_0 ? _GEN_636 : lvtReg_636; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1661 = io_wrEna_0 ? _GEN_637 : lvtReg_637; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1662 = io_wrEna_0 ? _GEN_638 : lvtReg_638; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1663 = io_wrEna_0 ? _GEN_639 : lvtReg_639; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1664 = io_wrEna_0 ? _GEN_640 : lvtReg_640; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1665 = io_wrEna_0 ? _GEN_641 : lvtReg_641; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1666 = io_wrEna_0 ? _GEN_642 : lvtReg_642; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1667 = io_wrEna_0 ? _GEN_643 : lvtReg_643; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1668 = io_wrEna_0 ? _GEN_644 : lvtReg_644; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1669 = io_wrEna_0 ? _GEN_645 : lvtReg_645; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1670 = io_wrEna_0 ? _GEN_646 : lvtReg_646; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1671 = io_wrEna_0 ? _GEN_647 : lvtReg_647; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1672 = io_wrEna_0 ? _GEN_648 : lvtReg_648; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1673 = io_wrEna_0 ? _GEN_649 : lvtReg_649; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1674 = io_wrEna_0 ? _GEN_650 : lvtReg_650; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1675 = io_wrEna_0 ? _GEN_651 : lvtReg_651; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1676 = io_wrEna_0 ? _GEN_652 : lvtReg_652; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1677 = io_wrEna_0 ? _GEN_653 : lvtReg_653; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1678 = io_wrEna_0 ? _GEN_654 : lvtReg_654; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1679 = io_wrEna_0 ? _GEN_655 : lvtReg_655; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1680 = io_wrEna_0 ? _GEN_656 : lvtReg_656; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1681 = io_wrEna_0 ? _GEN_657 : lvtReg_657; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1682 = io_wrEna_0 ? _GEN_658 : lvtReg_658; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1683 = io_wrEna_0 ? _GEN_659 : lvtReg_659; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1684 = io_wrEna_0 ? _GEN_660 : lvtReg_660; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1685 = io_wrEna_0 ? _GEN_661 : lvtReg_661; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1686 = io_wrEna_0 ? _GEN_662 : lvtReg_662; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1687 = io_wrEna_0 ? _GEN_663 : lvtReg_663; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1688 = io_wrEna_0 ? _GEN_664 : lvtReg_664; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1689 = io_wrEna_0 ? _GEN_665 : lvtReg_665; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1690 = io_wrEna_0 ? _GEN_666 : lvtReg_666; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1691 = io_wrEna_0 ? _GEN_667 : lvtReg_667; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1692 = io_wrEna_0 ? _GEN_668 : lvtReg_668; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1693 = io_wrEna_0 ? _GEN_669 : lvtReg_669; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1694 = io_wrEna_0 ? _GEN_670 : lvtReg_670; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1695 = io_wrEna_0 ? _GEN_671 : lvtReg_671; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1696 = io_wrEna_0 ? _GEN_672 : lvtReg_672; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1697 = io_wrEna_0 ? _GEN_673 : lvtReg_673; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1698 = io_wrEna_0 ? _GEN_674 : lvtReg_674; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1699 = io_wrEna_0 ? _GEN_675 : lvtReg_675; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1700 = io_wrEna_0 ? _GEN_676 : lvtReg_676; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1701 = io_wrEna_0 ? _GEN_677 : lvtReg_677; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1702 = io_wrEna_0 ? _GEN_678 : lvtReg_678; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1703 = io_wrEna_0 ? _GEN_679 : lvtReg_679; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1704 = io_wrEna_0 ? _GEN_680 : lvtReg_680; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1705 = io_wrEna_0 ? _GEN_681 : lvtReg_681; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1706 = io_wrEna_0 ? _GEN_682 : lvtReg_682; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1707 = io_wrEna_0 ? _GEN_683 : lvtReg_683; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1708 = io_wrEna_0 ? _GEN_684 : lvtReg_684; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1709 = io_wrEna_0 ? _GEN_685 : lvtReg_685; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1710 = io_wrEna_0 ? _GEN_686 : lvtReg_686; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1711 = io_wrEna_0 ? _GEN_687 : lvtReg_687; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1712 = io_wrEna_0 ? _GEN_688 : lvtReg_688; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1713 = io_wrEna_0 ? _GEN_689 : lvtReg_689; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1714 = io_wrEna_0 ? _GEN_690 : lvtReg_690; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1715 = io_wrEna_0 ? _GEN_691 : lvtReg_691; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1716 = io_wrEna_0 ? _GEN_692 : lvtReg_692; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1717 = io_wrEna_0 ? _GEN_693 : lvtReg_693; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1718 = io_wrEna_0 ? _GEN_694 : lvtReg_694; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1719 = io_wrEna_0 ? _GEN_695 : lvtReg_695; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1720 = io_wrEna_0 ? _GEN_696 : lvtReg_696; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1721 = io_wrEna_0 ? _GEN_697 : lvtReg_697; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1722 = io_wrEna_0 ? _GEN_698 : lvtReg_698; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1723 = io_wrEna_0 ? _GEN_699 : lvtReg_699; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1724 = io_wrEna_0 ? _GEN_700 : lvtReg_700; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1725 = io_wrEna_0 ? _GEN_701 : lvtReg_701; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1726 = io_wrEna_0 ? _GEN_702 : lvtReg_702; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1727 = io_wrEna_0 ? _GEN_703 : lvtReg_703; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1728 = io_wrEna_0 ? _GEN_704 : lvtReg_704; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1729 = io_wrEna_0 ? _GEN_705 : lvtReg_705; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1730 = io_wrEna_0 ? _GEN_706 : lvtReg_706; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1731 = io_wrEna_0 ? _GEN_707 : lvtReg_707; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1732 = io_wrEna_0 ? _GEN_708 : lvtReg_708; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1733 = io_wrEna_0 ? _GEN_709 : lvtReg_709; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1734 = io_wrEna_0 ? _GEN_710 : lvtReg_710; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1735 = io_wrEna_0 ? _GEN_711 : lvtReg_711; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1736 = io_wrEna_0 ? _GEN_712 : lvtReg_712; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1737 = io_wrEna_0 ? _GEN_713 : lvtReg_713; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1738 = io_wrEna_0 ? _GEN_714 : lvtReg_714; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1739 = io_wrEna_0 ? _GEN_715 : lvtReg_715; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1740 = io_wrEna_0 ? _GEN_716 : lvtReg_716; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1741 = io_wrEna_0 ? _GEN_717 : lvtReg_717; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1742 = io_wrEna_0 ? _GEN_718 : lvtReg_718; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1743 = io_wrEna_0 ? _GEN_719 : lvtReg_719; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1744 = io_wrEna_0 ? _GEN_720 : lvtReg_720; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1745 = io_wrEna_0 ? _GEN_721 : lvtReg_721; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1746 = io_wrEna_0 ? _GEN_722 : lvtReg_722; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1747 = io_wrEna_0 ? _GEN_723 : lvtReg_723; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1748 = io_wrEna_0 ? _GEN_724 : lvtReg_724; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1749 = io_wrEna_0 ? _GEN_725 : lvtReg_725; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1750 = io_wrEna_0 ? _GEN_726 : lvtReg_726; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1751 = io_wrEna_0 ? _GEN_727 : lvtReg_727; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1752 = io_wrEna_0 ? _GEN_728 : lvtReg_728; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1753 = io_wrEna_0 ? _GEN_729 : lvtReg_729; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1754 = io_wrEna_0 ? _GEN_730 : lvtReg_730; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1755 = io_wrEna_0 ? _GEN_731 : lvtReg_731; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1756 = io_wrEna_0 ? _GEN_732 : lvtReg_732; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1757 = io_wrEna_0 ? _GEN_733 : lvtReg_733; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1758 = io_wrEna_0 ? _GEN_734 : lvtReg_734; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1759 = io_wrEna_0 ? _GEN_735 : lvtReg_735; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1760 = io_wrEna_0 ? _GEN_736 : lvtReg_736; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1761 = io_wrEna_0 ? _GEN_737 : lvtReg_737; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1762 = io_wrEna_0 ? _GEN_738 : lvtReg_738; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1763 = io_wrEna_0 ? _GEN_739 : lvtReg_739; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1764 = io_wrEna_0 ? _GEN_740 : lvtReg_740; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1765 = io_wrEna_0 ? _GEN_741 : lvtReg_741; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1766 = io_wrEna_0 ? _GEN_742 : lvtReg_742; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1767 = io_wrEna_0 ? _GEN_743 : lvtReg_743; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1768 = io_wrEna_0 ? _GEN_744 : lvtReg_744; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1769 = io_wrEna_0 ? _GEN_745 : lvtReg_745; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1770 = io_wrEna_0 ? _GEN_746 : lvtReg_746; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1771 = io_wrEna_0 ? _GEN_747 : lvtReg_747; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1772 = io_wrEna_0 ? _GEN_748 : lvtReg_748; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1773 = io_wrEna_0 ? _GEN_749 : lvtReg_749; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1774 = io_wrEna_0 ? _GEN_750 : lvtReg_750; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1775 = io_wrEna_0 ? _GEN_751 : lvtReg_751; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1776 = io_wrEna_0 ? _GEN_752 : lvtReg_752; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1777 = io_wrEna_0 ? _GEN_753 : lvtReg_753; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1778 = io_wrEna_0 ? _GEN_754 : lvtReg_754; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1779 = io_wrEna_0 ? _GEN_755 : lvtReg_755; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1780 = io_wrEna_0 ? _GEN_756 : lvtReg_756; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1781 = io_wrEna_0 ? _GEN_757 : lvtReg_757; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1782 = io_wrEna_0 ? _GEN_758 : lvtReg_758; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1783 = io_wrEna_0 ? _GEN_759 : lvtReg_759; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1784 = io_wrEna_0 ? _GEN_760 : lvtReg_760; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1785 = io_wrEna_0 ? _GEN_761 : lvtReg_761; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1786 = io_wrEna_0 ? _GEN_762 : lvtReg_762; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1787 = io_wrEna_0 ? _GEN_763 : lvtReg_763; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1788 = io_wrEna_0 ? _GEN_764 : lvtReg_764; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1789 = io_wrEna_0 ? _GEN_765 : lvtReg_765; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1790 = io_wrEna_0 ? _GEN_766 : lvtReg_766; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1791 = io_wrEna_0 ? _GEN_767 : lvtReg_767; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1792 = io_wrEna_0 ? _GEN_768 : lvtReg_768; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1793 = io_wrEna_0 ? _GEN_769 : lvtReg_769; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1794 = io_wrEna_0 ? _GEN_770 : lvtReg_770; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1795 = io_wrEna_0 ? _GEN_771 : lvtReg_771; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1796 = io_wrEna_0 ? _GEN_772 : lvtReg_772; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1797 = io_wrEna_0 ? _GEN_773 : lvtReg_773; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1798 = io_wrEna_0 ? _GEN_774 : lvtReg_774; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1799 = io_wrEna_0 ? _GEN_775 : lvtReg_775; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1800 = io_wrEna_0 ? _GEN_776 : lvtReg_776; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1801 = io_wrEna_0 ? _GEN_777 : lvtReg_777; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1802 = io_wrEna_0 ? _GEN_778 : lvtReg_778; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1803 = io_wrEna_0 ? _GEN_779 : lvtReg_779; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1804 = io_wrEna_0 ? _GEN_780 : lvtReg_780; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1805 = io_wrEna_0 ? _GEN_781 : lvtReg_781; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1806 = io_wrEna_0 ? _GEN_782 : lvtReg_782; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1807 = io_wrEna_0 ? _GEN_783 : lvtReg_783; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1808 = io_wrEna_0 ? _GEN_784 : lvtReg_784; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1809 = io_wrEna_0 ? _GEN_785 : lvtReg_785; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1810 = io_wrEna_0 ? _GEN_786 : lvtReg_786; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1811 = io_wrEna_0 ? _GEN_787 : lvtReg_787; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1812 = io_wrEna_0 ? _GEN_788 : lvtReg_788; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1813 = io_wrEna_0 ? _GEN_789 : lvtReg_789; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1814 = io_wrEna_0 ? _GEN_790 : lvtReg_790; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1815 = io_wrEna_0 ? _GEN_791 : lvtReg_791; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1816 = io_wrEna_0 ? _GEN_792 : lvtReg_792; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1817 = io_wrEna_0 ? _GEN_793 : lvtReg_793; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1818 = io_wrEna_0 ? _GEN_794 : lvtReg_794; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1819 = io_wrEna_0 ? _GEN_795 : lvtReg_795; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1820 = io_wrEna_0 ? _GEN_796 : lvtReg_796; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1821 = io_wrEna_0 ? _GEN_797 : lvtReg_797; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1822 = io_wrEna_0 ? _GEN_798 : lvtReg_798; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1823 = io_wrEna_0 ? _GEN_799 : lvtReg_799; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1824 = io_wrEna_0 ? _GEN_800 : lvtReg_800; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1825 = io_wrEna_0 ? _GEN_801 : lvtReg_801; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1826 = io_wrEna_0 ? _GEN_802 : lvtReg_802; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1827 = io_wrEna_0 ? _GEN_803 : lvtReg_803; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1828 = io_wrEna_0 ? _GEN_804 : lvtReg_804; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1829 = io_wrEna_0 ? _GEN_805 : lvtReg_805; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1830 = io_wrEna_0 ? _GEN_806 : lvtReg_806; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1831 = io_wrEna_0 ? _GEN_807 : lvtReg_807; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1832 = io_wrEna_0 ? _GEN_808 : lvtReg_808; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1833 = io_wrEna_0 ? _GEN_809 : lvtReg_809; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1834 = io_wrEna_0 ? _GEN_810 : lvtReg_810; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1835 = io_wrEna_0 ? _GEN_811 : lvtReg_811; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1836 = io_wrEna_0 ? _GEN_812 : lvtReg_812; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1837 = io_wrEna_0 ? _GEN_813 : lvtReg_813; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1838 = io_wrEna_0 ? _GEN_814 : lvtReg_814; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1839 = io_wrEna_0 ? _GEN_815 : lvtReg_815; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1840 = io_wrEna_0 ? _GEN_816 : lvtReg_816; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1841 = io_wrEna_0 ? _GEN_817 : lvtReg_817; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1842 = io_wrEna_0 ? _GEN_818 : lvtReg_818; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1843 = io_wrEna_0 ? _GEN_819 : lvtReg_819; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1844 = io_wrEna_0 ? _GEN_820 : lvtReg_820; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1845 = io_wrEna_0 ? _GEN_821 : lvtReg_821; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1846 = io_wrEna_0 ? _GEN_822 : lvtReg_822; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1847 = io_wrEna_0 ? _GEN_823 : lvtReg_823; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1848 = io_wrEna_0 ? _GEN_824 : lvtReg_824; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1849 = io_wrEna_0 ? _GEN_825 : lvtReg_825; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1850 = io_wrEna_0 ? _GEN_826 : lvtReg_826; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1851 = io_wrEna_0 ? _GEN_827 : lvtReg_827; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1852 = io_wrEna_0 ? _GEN_828 : lvtReg_828; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1853 = io_wrEna_0 ? _GEN_829 : lvtReg_829; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1854 = io_wrEna_0 ? _GEN_830 : lvtReg_830; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1855 = io_wrEna_0 ? _GEN_831 : lvtReg_831; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1856 = io_wrEna_0 ? _GEN_832 : lvtReg_832; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1857 = io_wrEna_0 ? _GEN_833 : lvtReg_833; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1858 = io_wrEna_0 ? _GEN_834 : lvtReg_834; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1859 = io_wrEna_0 ? _GEN_835 : lvtReg_835; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1860 = io_wrEna_0 ? _GEN_836 : lvtReg_836; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1861 = io_wrEna_0 ? _GEN_837 : lvtReg_837; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1862 = io_wrEna_0 ? _GEN_838 : lvtReg_838; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1863 = io_wrEna_0 ? _GEN_839 : lvtReg_839; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1864 = io_wrEna_0 ? _GEN_840 : lvtReg_840; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1865 = io_wrEna_0 ? _GEN_841 : lvtReg_841; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1866 = io_wrEna_0 ? _GEN_842 : lvtReg_842; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1867 = io_wrEna_0 ? _GEN_843 : lvtReg_843; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1868 = io_wrEna_0 ? _GEN_844 : lvtReg_844; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1869 = io_wrEna_0 ? _GEN_845 : lvtReg_845; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1870 = io_wrEna_0 ? _GEN_846 : lvtReg_846; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1871 = io_wrEna_0 ? _GEN_847 : lvtReg_847; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1872 = io_wrEna_0 ? _GEN_848 : lvtReg_848; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1873 = io_wrEna_0 ? _GEN_849 : lvtReg_849; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1874 = io_wrEna_0 ? _GEN_850 : lvtReg_850; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1875 = io_wrEna_0 ? _GEN_851 : lvtReg_851; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1876 = io_wrEna_0 ? _GEN_852 : lvtReg_852; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1877 = io_wrEna_0 ? _GEN_853 : lvtReg_853; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1878 = io_wrEna_0 ? _GEN_854 : lvtReg_854; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1879 = io_wrEna_0 ? _GEN_855 : lvtReg_855; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1880 = io_wrEna_0 ? _GEN_856 : lvtReg_856; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1881 = io_wrEna_0 ? _GEN_857 : lvtReg_857; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1882 = io_wrEna_0 ? _GEN_858 : lvtReg_858; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1883 = io_wrEna_0 ? _GEN_859 : lvtReg_859; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1884 = io_wrEna_0 ? _GEN_860 : lvtReg_860; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1885 = io_wrEna_0 ? _GEN_861 : lvtReg_861; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1886 = io_wrEna_0 ? _GEN_862 : lvtReg_862; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1887 = io_wrEna_0 ? _GEN_863 : lvtReg_863; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1888 = io_wrEna_0 ? _GEN_864 : lvtReg_864; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1889 = io_wrEna_0 ? _GEN_865 : lvtReg_865; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1890 = io_wrEna_0 ? _GEN_866 : lvtReg_866; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1891 = io_wrEna_0 ? _GEN_867 : lvtReg_867; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1892 = io_wrEna_0 ? _GEN_868 : lvtReg_868; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1893 = io_wrEna_0 ? _GEN_869 : lvtReg_869; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1894 = io_wrEna_0 ? _GEN_870 : lvtReg_870; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1895 = io_wrEna_0 ? _GEN_871 : lvtReg_871; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1896 = io_wrEna_0 ? _GEN_872 : lvtReg_872; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1897 = io_wrEna_0 ? _GEN_873 : lvtReg_873; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1898 = io_wrEna_0 ? _GEN_874 : lvtReg_874; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1899 = io_wrEna_0 ? _GEN_875 : lvtReg_875; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1900 = io_wrEna_0 ? _GEN_876 : lvtReg_876; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1901 = io_wrEna_0 ? _GEN_877 : lvtReg_877; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1902 = io_wrEna_0 ? _GEN_878 : lvtReg_878; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1903 = io_wrEna_0 ? _GEN_879 : lvtReg_879; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1904 = io_wrEna_0 ? _GEN_880 : lvtReg_880; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1905 = io_wrEna_0 ? _GEN_881 : lvtReg_881; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1906 = io_wrEna_0 ? _GEN_882 : lvtReg_882; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1907 = io_wrEna_0 ? _GEN_883 : lvtReg_883; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1908 = io_wrEna_0 ? _GEN_884 : lvtReg_884; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1909 = io_wrEna_0 ? _GEN_885 : lvtReg_885; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1910 = io_wrEna_0 ? _GEN_886 : lvtReg_886; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1911 = io_wrEna_0 ? _GEN_887 : lvtReg_887; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1912 = io_wrEna_0 ? _GEN_888 : lvtReg_888; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1913 = io_wrEna_0 ? _GEN_889 : lvtReg_889; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1914 = io_wrEna_0 ? _GEN_890 : lvtReg_890; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1915 = io_wrEna_0 ? _GEN_891 : lvtReg_891; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1916 = io_wrEna_0 ? _GEN_892 : lvtReg_892; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1917 = io_wrEna_0 ? _GEN_893 : lvtReg_893; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1918 = io_wrEna_0 ? _GEN_894 : lvtReg_894; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1919 = io_wrEna_0 ? _GEN_895 : lvtReg_895; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1920 = io_wrEna_0 ? _GEN_896 : lvtReg_896; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1921 = io_wrEna_0 ? _GEN_897 : lvtReg_897; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1922 = io_wrEna_0 ? _GEN_898 : lvtReg_898; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1923 = io_wrEna_0 ? _GEN_899 : lvtReg_899; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1924 = io_wrEna_0 ? _GEN_900 : lvtReg_900; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1925 = io_wrEna_0 ? _GEN_901 : lvtReg_901; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1926 = io_wrEna_0 ? _GEN_902 : lvtReg_902; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1927 = io_wrEna_0 ? _GEN_903 : lvtReg_903; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1928 = io_wrEna_0 ? _GEN_904 : lvtReg_904; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1929 = io_wrEna_0 ? _GEN_905 : lvtReg_905; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1930 = io_wrEna_0 ? _GEN_906 : lvtReg_906; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1931 = io_wrEna_0 ? _GEN_907 : lvtReg_907; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1932 = io_wrEna_0 ? _GEN_908 : lvtReg_908; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1933 = io_wrEna_0 ? _GEN_909 : lvtReg_909; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1934 = io_wrEna_0 ? _GEN_910 : lvtReg_910; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1935 = io_wrEna_0 ? _GEN_911 : lvtReg_911; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1936 = io_wrEna_0 ? _GEN_912 : lvtReg_912; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1937 = io_wrEna_0 ? _GEN_913 : lvtReg_913; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1938 = io_wrEna_0 ? _GEN_914 : lvtReg_914; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1939 = io_wrEna_0 ? _GEN_915 : lvtReg_915; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1940 = io_wrEna_0 ? _GEN_916 : lvtReg_916; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1941 = io_wrEna_0 ? _GEN_917 : lvtReg_917; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1942 = io_wrEna_0 ? _GEN_918 : lvtReg_918; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1943 = io_wrEna_0 ? _GEN_919 : lvtReg_919; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1944 = io_wrEna_0 ? _GEN_920 : lvtReg_920; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1945 = io_wrEna_0 ? _GEN_921 : lvtReg_921; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1946 = io_wrEna_0 ? _GEN_922 : lvtReg_922; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1947 = io_wrEna_0 ? _GEN_923 : lvtReg_923; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1948 = io_wrEna_0 ? _GEN_924 : lvtReg_924; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1949 = io_wrEna_0 ? _GEN_925 : lvtReg_925; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1950 = io_wrEna_0 ? _GEN_926 : lvtReg_926; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1951 = io_wrEna_0 ? _GEN_927 : lvtReg_927; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1952 = io_wrEna_0 ? _GEN_928 : lvtReg_928; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1953 = io_wrEna_0 ? _GEN_929 : lvtReg_929; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1954 = io_wrEna_0 ? _GEN_930 : lvtReg_930; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1955 = io_wrEna_0 ? _GEN_931 : lvtReg_931; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1956 = io_wrEna_0 ? _GEN_932 : lvtReg_932; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1957 = io_wrEna_0 ? _GEN_933 : lvtReg_933; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1958 = io_wrEna_0 ? _GEN_934 : lvtReg_934; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1959 = io_wrEna_0 ? _GEN_935 : lvtReg_935; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1960 = io_wrEna_0 ? _GEN_936 : lvtReg_936; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1961 = io_wrEna_0 ? _GEN_937 : lvtReg_937; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1962 = io_wrEna_0 ? _GEN_938 : lvtReg_938; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1963 = io_wrEna_0 ? _GEN_939 : lvtReg_939; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1964 = io_wrEna_0 ? _GEN_940 : lvtReg_940; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1965 = io_wrEna_0 ? _GEN_941 : lvtReg_941; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1966 = io_wrEna_0 ? _GEN_942 : lvtReg_942; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1967 = io_wrEna_0 ? _GEN_943 : lvtReg_943; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1968 = io_wrEna_0 ? _GEN_944 : lvtReg_944; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1969 = io_wrEna_0 ? _GEN_945 : lvtReg_945; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1970 = io_wrEna_0 ? _GEN_946 : lvtReg_946; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1971 = io_wrEna_0 ? _GEN_947 : lvtReg_947; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1972 = io_wrEna_0 ? _GEN_948 : lvtReg_948; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1973 = io_wrEna_0 ? _GEN_949 : lvtReg_949; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1974 = io_wrEna_0 ? _GEN_950 : lvtReg_950; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1975 = io_wrEna_0 ? _GEN_951 : lvtReg_951; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1976 = io_wrEna_0 ? _GEN_952 : lvtReg_952; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1977 = io_wrEna_0 ? _GEN_953 : lvtReg_953; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1978 = io_wrEna_0 ? _GEN_954 : lvtReg_954; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1979 = io_wrEna_0 ? _GEN_955 : lvtReg_955; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1980 = io_wrEna_0 ? _GEN_956 : lvtReg_956; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1981 = io_wrEna_0 ? _GEN_957 : lvtReg_957; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1982 = io_wrEna_0 ? _GEN_958 : lvtReg_958; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1983 = io_wrEna_0 ? _GEN_959 : lvtReg_959; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1984 = io_wrEna_0 ? _GEN_960 : lvtReg_960; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1985 = io_wrEna_0 ? _GEN_961 : lvtReg_961; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1986 = io_wrEna_0 ? _GEN_962 : lvtReg_962; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1987 = io_wrEna_0 ? _GEN_963 : lvtReg_963; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1988 = io_wrEna_0 ? _GEN_964 : lvtReg_964; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1989 = io_wrEna_0 ? _GEN_965 : lvtReg_965; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1990 = io_wrEna_0 ? _GEN_966 : lvtReg_966; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1991 = io_wrEna_0 ? _GEN_967 : lvtReg_967; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1992 = io_wrEna_0 ? _GEN_968 : lvtReg_968; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1993 = io_wrEna_0 ? _GEN_969 : lvtReg_969; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1994 = io_wrEna_0 ? _GEN_970 : lvtReg_970; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1995 = io_wrEna_0 ? _GEN_971 : lvtReg_971; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1996 = io_wrEna_0 ? _GEN_972 : lvtReg_972; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1997 = io_wrEna_0 ? _GEN_973 : lvtReg_973; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1998 = io_wrEna_0 ? _GEN_974 : lvtReg_974; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1999 = io_wrEna_0 ? _GEN_975 : lvtReg_975; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2000 = io_wrEna_0 ? _GEN_976 : lvtReg_976; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2001 = io_wrEna_0 ? _GEN_977 : lvtReg_977; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2002 = io_wrEna_0 ? _GEN_978 : lvtReg_978; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2003 = io_wrEna_0 ? _GEN_979 : lvtReg_979; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2004 = io_wrEna_0 ? _GEN_980 : lvtReg_980; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2005 = io_wrEna_0 ? _GEN_981 : lvtReg_981; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2006 = io_wrEna_0 ? _GEN_982 : lvtReg_982; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2007 = io_wrEna_0 ? _GEN_983 : lvtReg_983; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2008 = io_wrEna_0 ? _GEN_984 : lvtReg_984; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2009 = io_wrEna_0 ? _GEN_985 : lvtReg_985; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2010 = io_wrEna_0 ? _GEN_986 : lvtReg_986; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2011 = io_wrEna_0 ? _GEN_987 : lvtReg_987; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2012 = io_wrEna_0 ? _GEN_988 : lvtReg_988; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2013 = io_wrEna_0 ? _GEN_989 : lvtReg_989; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2014 = io_wrEna_0 ? _GEN_990 : lvtReg_990; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2015 = io_wrEna_0 ? _GEN_991 : lvtReg_991; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2016 = io_wrEna_0 ? _GEN_992 : lvtReg_992; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2017 = io_wrEna_0 ? _GEN_993 : lvtReg_993; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2018 = io_wrEna_0 ? _GEN_994 : lvtReg_994; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2019 = io_wrEna_0 ? _GEN_995 : lvtReg_995; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2020 = io_wrEna_0 ? _GEN_996 : lvtReg_996; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2021 = io_wrEna_0 ? _GEN_997 : lvtReg_997; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2022 = io_wrEna_0 ? _GEN_998 : lvtReg_998; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2023 = io_wrEna_0 ? _GEN_999 : lvtReg_999; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2024 = io_wrEna_0 ? _GEN_1000 : lvtReg_1000; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2025 = io_wrEna_0 ? _GEN_1001 : lvtReg_1001; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2026 = io_wrEna_0 ? _GEN_1002 : lvtReg_1002; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2027 = io_wrEna_0 ? _GEN_1003 : lvtReg_1003; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2028 = io_wrEna_0 ? _GEN_1004 : lvtReg_1004; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2029 = io_wrEna_0 ? _GEN_1005 : lvtReg_1005; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2030 = io_wrEna_0 ? _GEN_1006 : lvtReg_1006; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2031 = io_wrEna_0 ? _GEN_1007 : lvtReg_1007; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2032 = io_wrEna_0 ? _GEN_1008 : lvtReg_1008; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2033 = io_wrEna_0 ? _GEN_1009 : lvtReg_1009; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2034 = io_wrEna_0 ? _GEN_1010 : lvtReg_1010; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2035 = io_wrEna_0 ? _GEN_1011 : lvtReg_1011; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2036 = io_wrEna_0 ? _GEN_1012 : lvtReg_1012; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2037 = io_wrEna_0 ? _GEN_1013 : lvtReg_1013; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2038 = io_wrEna_0 ? _GEN_1014 : lvtReg_1014; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2039 = io_wrEna_0 ? _GEN_1015 : lvtReg_1015; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2040 = io_wrEna_0 ? _GEN_1016 : lvtReg_1016; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2041 = io_wrEna_0 ? _GEN_1017 : lvtReg_1017; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2042 = io_wrEna_0 ? _GEN_1018 : lvtReg_1018; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2043 = io_wrEna_0 ? _GEN_1019 : lvtReg_1019; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2044 = io_wrEna_0 ? _GEN_1020 : lvtReg_1020; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2045 = io_wrEna_0 ? _GEN_1021 : lvtReg_1021; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2046 = io_wrEna_0 ? _GEN_1022 : lvtReg_1022; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2047 = io_wrEna_0 ? _GEN_1023 : lvtReg_1023; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_4097 = 10'h1 == io_rdAddr_0 ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4098 = 10'h2 == io_rdAddr_0 ? lvtReg_2 : _GEN_4097; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4099 = 10'h3 == io_rdAddr_0 ? lvtReg_3 : _GEN_4098; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4100 = 10'h4 == io_rdAddr_0 ? lvtReg_4 : _GEN_4099; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4101 = 10'h5 == io_rdAddr_0 ? lvtReg_5 : _GEN_4100; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4102 = 10'h6 == io_rdAddr_0 ? lvtReg_6 : _GEN_4101; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4103 = 10'h7 == io_rdAddr_0 ? lvtReg_7 : _GEN_4102; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4104 = 10'h8 == io_rdAddr_0 ? lvtReg_8 : _GEN_4103; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4105 = 10'h9 == io_rdAddr_0 ? lvtReg_9 : _GEN_4104; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4106 = 10'ha == io_rdAddr_0 ? lvtReg_10 : _GEN_4105; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4107 = 10'hb == io_rdAddr_0 ? lvtReg_11 : _GEN_4106; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4108 = 10'hc == io_rdAddr_0 ? lvtReg_12 : _GEN_4107; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4109 = 10'hd == io_rdAddr_0 ? lvtReg_13 : _GEN_4108; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4110 = 10'he == io_rdAddr_0 ? lvtReg_14 : _GEN_4109; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4111 = 10'hf == io_rdAddr_0 ? lvtReg_15 : _GEN_4110; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4112 = 10'h10 == io_rdAddr_0 ? lvtReg_16 : _GEN_4111; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4113 = 10'h11 == io_rdAddr_0 ? lvtReg_17 : _GEN_4112; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4114 = 10'h12 == io_rdAddr_0 ? lvtReg_18 : _GEN_4113; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4115 = 10'h13 == io_rdAddr_0 ? lvtReg_19 : _GEN_4114; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4116 = 10'h14 == io_rdAddr_0 ? lvtReg_20 : _GEN_4115; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4117 = 10'h15 == io_rdAddr_0 ? lvtReg_21 : _GEN_4116; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4118 = 10'h16 == io_rdAddr_0 ? lvtReg_22 : _GEN_4117; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4119 = 10'h17 == io_rdAddr_0 ? lvtReg_23 : _GEN_4118; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4120 = 10'h18 == io_rdAddr_0 ? lvtReg_24 : _GEN_4119; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4121 = 10'h19 == io_rdAddr_0 ? lvtReg_25 : _GEN_4120; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4122 = 10'h1a == io_rdAddr_0 ? lvtReg_26 : _GEN_4121; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4123 = 10'h1b == io_rdAddr_0 ? lvtReg_27 : _GEN_4122; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4124 = 10'h1c == io_rdAddr_0 ? lvtReg_28 : _GEN_4123; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4125 = 10'h1d == io_rdAddr_0 ? lvtReg_29 : _GEN_4124; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4126 = 10'h1e == io_rdAddr_0 ? lvtReg_30 : _GEN_4125; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4127 = 10'h1f == io_rdAddr_0 ? lvtReg_31 : _GEN_4126; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4128 = 10'h20 == io_rdAddr_0 ? lvtReg_32 : _GEN_4127; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4129 = 10'h21 == io_rdAddr_0 ? lvtReg_33 : _GEN_4128; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4130 = 10'h22 == io_rdAddr_0 ? lvtReg_34 : _GEN_4129; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4131 = 10'h23 == io_rdAddr_0 ? lvtReg_35 : _GEN_4130; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4132 = 10'h24 == io_rdAddr_0 ? lvtReg_36 : _GEN_4131; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4133 = 10'h25 == io_rdAddr_0 ? lvtReg_37 : _GEN_4132; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4134 = 10'h26 == io_rdAddr_0 ? lvtReg_38 : _GEN_4133; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4135 = 10'h27 == io_rdAddr_0 ? lvtReg_39 : _GEN_4134; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4136 = 10'h28 == io_rdAddr_0 ? lvtReg_40 : _GEN_4135; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4137 = 10'h29 == io_rdAddr_0 ? lvtReg_41 : _GEN_4136; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4138 = 10'h2a == io_rdAddr_0 ? lvtReg_42 : _GEN_4137; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4139 = 10'h2b == io_rdAddr_0 ? lvtReg_43 : _GEN_4138; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4140 = 10'h2c == io_rdAddr_0 ? lvtReg_44 : _GEN_4139; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4141 = 10'h2d == io_rdAddr_0 ? lvtReg_45 : _GEN_4140; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4142 = 10'h2e == io_rdAddr_0 ? lvtReg_46 : _GEN_4141; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4143 = 10'h2f == io_rdAddr_0 ? lvtReg_47 : _GEN_4142; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4144 = 10'h30 == io_rdAddr_0 ? lvtReg_48 : _GEN_4143; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4145 = 10'h31 == io_rdAddr_0 ? lvtReg_49 : _GEN_4144; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4146 = 10'h32 == io_rdAddr_0 ? lvtReg_50 : _GEN_4145; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4147 = 10'h33 == io_rdAddr_0 ? lvtReg_51 : _GEN_4146; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4148 = 10'h34 == io_rdAddr_0 ? lvtReg_52 : _GEN_4147; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4149 = 10'h35 == io_rdAddr_0 ? lvtReg_53 : _GEN_4148; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4150 = 10'h36 == io_rdAddr_0 ? lvtReg_54 : _GEN_4149; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4151 = 10'h37 == io_rdAddr_0 ? lvtReg_55 : _GEN_4150; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4152 = 10'h38 == io_rdAddr_0 ? lvtReg_56 : _GEN_4151; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4153 = 10'h39 == io_rdAddr_0 ? lvtReg_57 : _GEN_4152; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4154 = 10'h3a == io_rdAddr_0 ? lvtReg_58 : _GEN_4153; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4155 = 10'h3b == io_rdAddr_0 ? lvtReg_59 : _GEN_4154; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4156 = 10'h3c == io_rdAddr_0 ? lvtReg_60 : _GEN_4155; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4157 = 10'h3d == io_rdAddr_0 ? lvtReg_61 : _GEN_4156; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4158 = 10'h3e == io_rdAddr_0 ? lvtReg_62 : _GEN_4157; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4159 = 10'h3f == io_rdAddr_0 ? lvtReg_63 : _GEN_4158; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4160 = 10'h40 == io_rdAddr_0 ? lvtReg_64 : _GEN_4159; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4161 = 10'h41 == io_rdAddr_0 ? lvtReg_65 : _GEN_4160; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4162 = 10'h42 == io_rdAddr_0 ? lvtReg_66 : _GEN_4161; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4163 = 10'h43 == io_rdAddr_0 ? lvtReg_67 : _GEN_4162; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4164 = 10'h44 == io_rdAddr_0 ? lvtReg_68 : _GEN_4163; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4165 = 10'h45 == io_rdAddr_0 ? lvtReg_69 : _GEN_4164; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4166 = 10'h46 == io_rdAddr_0 ? lvtReg_70 : _GEN_4165; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4167 = 10'h47 == io_rdAddr_0 ? lvtReg_71 : _GEN_4166; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4168 = 10'h48 == io_rdAddr_0 ? lvtReg_72 : _GEN_4167; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4169 = 10'h49 == io_rdAddr_0 ? lvtReg_73 : _GEN_4168; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4170 = 10'h4a == io_rdAddr_0 ? lvtReg_74 : _GEN_4169; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4171 = 10'h4b == io_rdAddr_0 ? lvtReg_75 : _GEN_4170; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4172 = 10'h4c == io_rdAddr_0 ? lvtReg_76 : _GEN_4171; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4173 = 10'h4d == io_rdAddr_0 ? lvtReg_77 : _GEN_4172; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4174 = 10'h4e == io_rdAddr_0 ? lvtReg_78 : _GEN_4173; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4175 = 10'h4f == io_rdAddr_0 ? lvtReg_79 : _GEN_4174; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4176 = 10'h50 == io_rdAddr_0 ? lvtReg_80 : _GEN_4175; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4177 = 10'h51 == io_rdAddr_0 ? lvtReg_81 : _GEN_4176; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4178 = 10'h52 == io_rdAddr_0 ? lvtReg_82 : _GEN_4177; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4179 = 10'h53 == io_rdAddr_0 ? lvtReg_83 : _GEN_4178; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4180 = 10'h54 == io_rdAddr_0 ? lvtReg_84 : _GEN_4179; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4181 = 10'h55 == io_rdAddr_0 ? lvtReg_85 : _GEN_4180; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4182 = 10'h56 == io_rdAddr_0 ? lvtReg_86 : _GEN_4181; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4183 = 10'h57 == io_rdAddr_0 ? lvtReg_87 : _GEN_4182; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4184 = 10'h58 == io_rdAddr_0 ? lvtReg_88 : _GEN_4183; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4185 = 10'h59 == io_rdAddr_0 ? lvtReg_89 : _GEN_4184; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4186 = 10'h5a == io_rdAddr_0 ? lvtReg_90 : _GEN_4185; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4187 = 10'h5b == io_rdAddr_0 ? lvtReg_91 : _GEN_4186; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4188 = 10'h5c == io_rdAddr_0 ? lvtReg_92 : _GEN_4187; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4189 = 10'h5d == io_rdAddr_0 ? lvtReg_93 : _GEN_4188; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4190 = 10'h5e == io_rdAddr_0 ? lvtReg_94 : _GEN_4189; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4191 = 10'h5f == io_rdAddr_0 ? lvtReg_95 : _GEN_4190; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4192 = 10'h60 == io_rdAddr_0 ? lvtReg_96 : _GEN_4191; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4193 = 10'h61 == io_rdAddr_0 ? lvtReg_97 : _GEN_4192; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4194 = 10'h62 == io_rdAddr_0 ? lvtReg_98 : _GEN_4193; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4195 = 10'h63 == io_rdAddr_0 ? lvtReg_99 : _GEN_4194; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4196 = 10'h64 == io_rdAddr_0 ? lvtReg_100 : _GEN_4195; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4197 = 10'h65 == io_rdAddr_0 ? lvtReg_101 : _GEN_4196; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4198 = 10'h66 == io_rdAddr_0 ? lvtReg_102 : _GEN_4197; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4199 = 10'h67 == io_rdAddr_0 ? lvtReg_103 : _GEN_4198; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4200 = 10'h68 == io_rdAddr_0 ? lvtReg_104 : _GEN_4199; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4201 = 10'h69 == io_rdAddr_0 ? lvtReg_105 : _GEN_4200; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4202 = 10'h6a == io_rdAddr_0 ? lvtReg_106 : _GEN_4201; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4203 = 10'h6b == io_rdAddr_0 ? lvtReg_107 : _GEN_4202; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4204 = 10'h6c == io_rdAddr_0 ? lvtReg_108 : _GEN_4203; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4205 = 10'h6d == io_rdAddr_0 ? lvtReg_109 : _GEN_4204; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4206 = 10'h6e == io_rdAddr_0 ? lvtReg_110 : _GEN_4205; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4207 = 10'h6f == io_rdAddr_0 ? lvtReg_111 : _GEN_4206; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4208 = 10'h70 == io_rdAddr_0 ? lvtReg_112 : _GEN_4207; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4209 = 10'h71 == io_rdAddr_0 ? lvtReg_113 : _GEN_4208; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4210 = 10'h72 == io_rdAddr_0 ? lvtReg_114 : _GEN_4209; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4211 = 10'h73 == io_rdAddr_0 ? lvtReg_115 : _GEN_4210; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4212 = 10'h74 == io_rdAddr_0 ? lvtReg_116 : _GEN_4211; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4213 = 10'h75 == io_rdAddr_0 ? lvtReg_117 : _GEN_4212; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4214 = 10'h76 == io_rdAddr_0 ? lvtReg_118 : _GEN_4213; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4215 = 10'h77 == io_rdAddr_0 ? lvtReg_119 : _GEN_4214; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4216 = 10'h78 == io_rdAddr_0 ? lvtReg_120 : _GEN_4215; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4217 = 10'h79 == io_rdAddr_0 ? lvtReg_121 : _GEN_4216; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4218 = 10'h7a == io_rdAddr_0 ? lvtReg_122 : _GEN_4217; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4219 = 10'h7b == io_rdAddr_0 ? lvtReg_123 : _GEN_4218; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4220 = 10'h7c == io_rdAddr_0 ? lvtReg_124 : _GEN_4219; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4221 = 10'h7d == io_rdAddr_0 ? lvtReg_125 : _GEN_4220; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4222 = 10'h7e == io_rdAddr_0 ? lvtReg_126 : _GEN_4221; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4223 = 10'h7f == io_rdAddr_0 ? lvtReg_127 : _GEN_4222; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4224 = 10'h80 == io_rdAddr_0 ? lvtReg_128 : _GEN_4223; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4225 = 10'h81 == io_rdAddr_0 ? lvtReg_129 : _GEN_4224; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4226 = 10'h82 == io_rdAddr_0 ? lvtReg_130 : _GEN_4225; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4227 = 10'h83 == io_rdAddr_0 ? lvtReg_131 : _GEN_4226; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4228 = 10'h84 == io_rdAddr_0 ? lvtReg_132 : _GEN_4227; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4229 = 10'h85 == io_rdAddr_0 ? lvtReg_133 : _GEN_4228; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4230 = 10'h86 == io_rdAddr_0 ? lvtReg_134 : _GEN_4229; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4231 = 10'h87 == io_rdAddr_0 ? lvtReg_135 : _GEN_4230; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4232 = 10'h88 == io_rdAddr_0 ? lvtReg_136 : _GEN_4231; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4233 = 10'h89 == io_rdAddr_0 ? lvtReg_137 : _GEN_4232; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4234 = 10'h8a == io_rdAddr_0 ? lvtReg_138 : _GEN_4233; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4235 = 10'h8b == io_rdAddr_0 ? lvtReg_139 : _GEN_4234; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4236 = 10'h8c == io_rdAddr_0 ? lvtReg_140 : _GEN_4235; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4237 = 10'h8d == io_rdAddr_0 ? lvtReg_141 : _GEN_4236; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4238 = 10'h8e == io_rdAddr_0 ? lvtReg_142 : _GEN_4237; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4239 = 10'h8f == io_rdAddr_0 ? lvtReg_143 : _GEN_4238; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4240 = 10'h90 == io_rdAddr_0 ? lvtReg_144 : _GEN_4239; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4241 = 10'h91 == io_rdAddr_0 ? lvtReg_145 : _GEN_4240; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4242 = 10'h92 == io_rdAddr_0 ? lvtReg_146 : _GEN_4241; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4243 = 10'h93 == io_rdAddr_0 ? lvtReg_147 : _GEN_4242; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4244 = 10'h94 == io_rdAddr_0 ? lvtReg_148 : _GEN_4243; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4245 = 10'h95 == io_rdAddr_0 ? lvtReg_149 : _GEN_4244; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4246 = 10'h96 == io_rdAddr_0 ? lvtReg_150 : _GEN_4245; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4247 = 10'h97 == io_rdAddr_0 ? lvtReg_151 : _GEN_4246; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4248 = 10'h98 == io_rdAddr_0 ? lvtReg_152 : _GEN_4247; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4249 = 10'h99 == io_rdAddr_0 ? lvtReg_153 : _GEN_4248; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4250 = 10'h9a == io_rdAddr_0 ? lvtReg_154 : _GEN_4249; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4251 = 10'h9b == io_rdAddr_0 ? lvtReg_155 : _GEN_4250; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4252 = 10'h9c == io_rdAddr_0 ? lvtReg_156 : _GEN_4251; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4253 = 10'h9d == io_rdAddr_0 ? lvtReg_157 : _GEN_4252; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4254 = 10'h9e == io_rdAddr_0 ? lvtReg_158 : _GEN_4253; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4255 = 10'h9f == io_rdAddr_0 ? lvtReg_159 : _GEN_4254; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4256 = 10'ha0 == io_rdAddr_0 ? lvtReg_160 : _GEN_4255; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4257 = 10'ha1 == io_rdAddr_0 ? lvtReg_161 : _GEN_4256; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4258 = 10'ha2 == io_rdAddr_0 ? lvtReg_162 : _GEN_4257; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4259 = 10'ha3 == io_rdAddr_0 ? lvtReg_163 : _GEN_4258; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4260 = 10'ha4 == io_rdAddr_0 ? lvtReg_164 : _GEN_4259; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4261 = 10'ha5 == io_rdAddr_0 ? lvtReg_165 : _GEN_4260; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4262 = 10'ha6 == io_rdAddr_0 ? lvtReg_166 : _GEN_4261; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4263 = 10'ha7 == io_rdAddr_0 ? lvtReg_167 : _GEN_4262; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4264 = 10'ha8 == io_rdAddr_0 ? lvtReg_168 : _GEN_4263; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4265 = 10'ha9 == io_rdAddr_0 ? lvtReg_169 : _GEN_4264; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4266 = 10'haa == io_rdAddr_0 ? lvtReg_170 : _GEN_4265; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4267 = 10'hab == io_rdAddr_0 ? lvtReg_171 : _GEN_4266; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4268 = 10'hac == io_rdAddr_0 ? lvtReg_172 : _GEN_4267; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4269 = 10'had == io_rdAddr_0 ? lvtReg_173 : _GEN_4268; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4270 = 10'hae == io_rdAddr_0 ? lvtReg_174 : _GEN_4269; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4271 = 10'haf == io_rdAddr_0 ? lvtReg_175 : _GEN_4270; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4272 = 10'hb0 == io_rdAddr_0 ? lvtReg_176 : _GEN_4271; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4273 = 10'hb1 == io_rdAddr_0 ? lvtReg_177 : _GEN_4272; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4274 = 10'hb2 == io_rdAddr_0 ? lvtReg_178 : _GEN_4273; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4275 = 10'hb3 == io_rdAddr_0 ? lvtReg_179 : _GEN_4274; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4276 = 10'hb4 == io_rdAddr_0 ? lvtReg_180 : _GEN_4275; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4277 = 10'hb5 == io_rdAddr_0 ? lvtReg_181 : _GEN_4276; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4278 = 10'hb6 == io_rdAddr_0 ? lvtReg_182 : _GEN_4277; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4279 = 10'hb7 == io_rdAddr_0 ? lvtReg_183 : _GEN_4278; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4280 = 10'hb8 == io_rdAddr_0 ? lvtReg_184 : _GEN_4279; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4281 = 10'hb9 == io_rdAddr_0 ? lvtReg_185 : _GEN_4280; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4282 = 10'hba == io_rdAddr_0 ? lvtReg_186 : _GEN_4281; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4283 = 10'hbb == io_rdAddr_0 ? lvtReg_187 : _GEN_4282; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4284 = 10'hbc == io_rdAddr_0 ? lvtReg_188 : _GEN_4283; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4285 = 10'hbd == io_rdAddr_0 ? lvtReg_189 : _GEN_4284; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4286 = 10'hbe == io_rdAddr_0 ? lvtReg_190 : _GEN_4285; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4287 = 10'hbf == io_rdAddr_0 ? lvtReg_191 : _GEN_4286; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4288 = 10'hc0 == io_rdAddr_0 ? lvtReg_192 : _GEN_4287; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4289 = 10'hc1 == io_rdAddr_0 ? lvtReg_193 : _GEN_4288; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4290 = 10'hc2 == io_rdAddr_0 ? lvtReg_194 : _GEN_4289; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4291 = 10'hc3 == io_rdAddr_0 ? lvtReg_195 : _GEN_4290; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4292 = 10'hc4 == io_rdAddr_0 ? lvtReg_196 : _GEN_4291; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4293 = 10'hc5 == io_rdAddr_0 ? lvtReg_197 : _GEN_4292; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4294 = 10'hc6 == io_rdAddr_0 ? lvtReg_198 : _GEN_4293; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4295 = 10'hc7 == io_rdAddr_0 ? lvtReg_199 : _GEN_4294; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4296 = 10'hc8 == io_rdAddr_0 ? lvtReg_200 : _GEN_4295; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4297 = 10'hc9 == io_rdAddr_0 ? lvtReg_201 : _GEN_4296; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4298 = 10'hca == io_rdAddr_0 ? lvtReg_202 : _GEN_4297; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4299 = 10'hcb == io_rdAddr_0 ? lvtReg_203 : _GEN_4298; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4300 = 10'hcc == io_rdAddr_0 ? lvtReg_204 : _GEN_4299; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4301 = 10'hcd == io_rdAddr_0 ? lvtReg_205 : _GEN_4300; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4302 = 10'hce == io_rdAddr_0 ? lvtReg_206 : _GEN_4301; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4303 = 10'hcf == io_rdAddr_0 ? lvtReg_207 : _GEN_4302; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4304 = 10'hd0 == io_rdAddr_0 ? lvtReg_208 : _GEN_4303; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4305 = 10'hd1 == io_rdAddr_0 ? lvtReg_209 : _GEN_4304; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4306 = 10'hd2 == io_rdAddr_0 ? lvtReg_210 : _GEN_4305; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4307 = 10'hd3 == io_rdAddr_0 ? lvtReg_211 : _GEN_4306; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4308 = 10'hd4 == io_rdAddr_0 ? lvtReg_212 : _GEN_4307; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4309 = 10'hd5 == io_rdAddr_0 ? lvtReg_213 : _GEN_4308; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4310 = 10'hd6 == io_rdAddr_0 ? lvtReg_214 : _GEN_4309; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4311 = 10'hd7 == io_rdAddr_0 ? lvtReg_215 : _GEN_4310; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4312 = 10'hd8 == io_rdAddr_0 ? lvtReg_216 : _GEN_4311; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4313 = 10'hd9 == io_rdAddr_0 ? lvtReg_217 : _GEN_4312; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4314 = 10'hda == io_rdAddr_0 ? lvtReg_218 : _GEN_4313; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4315 = 10'hdb == io_rdAddr_0 ? lvtReg_219 : _GEN_4314; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4316 = 10'hdc == io_rdAddr_0 ? lvtReg_220 : _GEN_4315; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4317 = 10'hdd == io_rdAddr_0 ? lvtReg_221 : _GEN_4316; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4318 = 10'hde == io_rdAddr_0 ? lvtReg_222 : _GEN_4317; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4319 = 10'hdf == io_rdAddr_0 ? lvtReg_223 : _GEN_4318; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4320 = 10'he0 == io_rdAddr_0 ? lvtReg_224 : _GEN_4319; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4321 = 10'he1 == io_rdAddr_0 ? lvtReg_225 : _GEN_4320; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4322 = 10'he2 == io_rdAddr_0 ? lvtReg_226 : _GEN_4321; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4323 = 10'he3 == io_rdAddr_0 ? lvtReg_227 : _GEN_4322; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4324 = 10'he4 == io_rdAddr_0 ? lvtReg_228 : _GEN_4323; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4325 = 10'he5 == io_rdAddr_0 ? lvtReg_229 : _GEN_4324; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4326 = 10'he6 == io_rdAddr_0 ? lvtReg_230 : _GEN_4325; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4327 = 10'he7 == io_rdAddr_0 ? lvtReg_231 : _GEN_4326; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4328 = 10'he8 == io_rdAddr_0 ? lvtReg_232 : _GEN_4327; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4329 = 10'he9 == io_rdAddr_0 ? lvtReg_233 : _GEN_4328; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4330 = 10'hea == io_rdAddr_0 ? lvtReg_234 : _GEN_4329; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4331 = 10'heb == io_rdAddr_0 ? lvtReg_235 : _GEN_4330; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4332 = 10'hec == io_rdAddr_0 ? lvtReg_236 : _GEN_4331; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4333 = 10'hed == io_rdAddr_0 ? lvtReg_237 : _GEN_4332; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4334 = 10'hee == io_rdAddr_0 ? lvtReg_238 : _GEN_4333; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4335 = 10'hef == io_rdAddr_0 ? lvtReg_239 : _GEN_4334; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4336 = 10'hf0 == io_rdAddr_0 ? lvtReg_240 : _GEN_4335; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4337 = 10'hf1 == io_rdAddr_0 ? lvtReg_241 : _GEN_4336; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4338 = 10'hf2 == io_rdAddr_0 ? lvtReg_242 : _GEN_4337; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4339 = 10'hf3 == io_rdAddr_0 ? lvtReg_243 : _GEN_4338; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4340 = 10'hf4 == io_rdAddr_0 ? lvtReg_244 : _GEN_4339; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4341 = 10'hf5 == io_rdAddr_0 ? lvtReg_245 : _GEN_4340; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4342 = 10'hf6 == io_rdAddr_0 ? lvtReg_246 : _GEN_4341; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4343 = 10'hf7 == io_rdAddr_0 ? lvtReg_247 : _GEN_4342; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4344 = 10'hf8 == io_rdAddr_0 ? lvtReg_248 : _GEN_4343; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4345 = 10'hf9 == io_rdAddr_0 ? lvtReg_249 : _GEN_4344; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4346 = 10'hfa == io_rdAddr_0 ? lvtReg_250 : _GEN_4345; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4347 = 10'hfb == io_rdAddr_0 ? lvtReg_251 : _GEN_4346; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4348 = 10'hfc == io_rdAddr_0 ? lvtReg_252 : _GEN_4347; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4349 = 10'hfd == io_rdAddr_0 ? lvtReg_253 : _GEN_4348; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4350 = 10'hfe == io_rdAddr_0 ? lvtReg_254 : _GEN_4349; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4351 = 10'hff == io_rdAddr_0 ? lvtReg_255 : _GEN_4350; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4352 = 10'h100 == io_rdAddr_0 ? lvtReg_256 : _GEN_4351; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4353 = 10'h101 == io_rdAddr_0 ? lvtReg_257 : _GEN_4352; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4354 = 10'h102 == io_rdAddr_0 ? lvtReg_258 : _GEN_4353; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4355 = 10'h103 == io_rdAddr_0 ? lvtReg_259 : _GEN_4354; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4356 = 10'h104 == io_rdAddr_0 ? lvtReg_260 : _GEN_4355; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4357 = 10'h105 == io_rdAddr_0 ? lvtReg_261 : _GEN_4356; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4358 = 10'h106 == io_rdAddr_0 ? lvtReg_262 : _GEN_4357; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4359 = 10'h107 == io_rdAddr_0 ? lvtReg_263 : _GEN_4358; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4360 = 10'h108 == io_rdAddr_0 ? lvtReg_264 : _GEN_4359; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4361 = 10'h109 == io_rdAddr_0 ? lvtReg_265 : _GEN_4360; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4362 = 10'h10a == io_rdAddr_0 ? lvtReg_266 : _GEN_4361; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4363 = 10'h10b == io_rdAddr_0 ? lvtReg_267 : _GEN_4362; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4364 = 10'h10c == io_rdAddr_0 ? lvtReg_268 : _GEN_4363; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4365 = 10'h10d == io_rdAddr_0 ? lvtReg_269 : _GEN_4364; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4366 = 10'h10e == io_rdAddr_0 ? lvtReg_270 : _GEN_4365; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4367 = 10'h10f == io_rdAddr_0 ? lvtReg_271 : _GEN_4366; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4368 = 10'h110 == io_rdAddr_0 ? lvtReg_272 : _GEN_4367; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4369 = 10'h111 == io_rdAddr_0 ? lvtReg_273 : _GEN_4368; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4370 = 10'h112 == io_rdAddr_0 ? lvtReg_274 : _GEN_4369; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4371 = 10'h113 == io_rdAddr_0 ? lvtReg_275 : _GEN_4370; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4372 = 10'h114 == io_rdAddr_0 ? lvtReg_276 : _GEN_4371; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4373 = 10'h115 == io_rdAddr_0 ? lvtReg_277 : _GEN_4372; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4374 = 10'h116 == io_rdAddr_0 ? lvtReg_278 : _GEN_4373; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4375 = 10'h117 == io_rdAddr_0 ? lvtReg_279 : _GEN_4374; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4376 = 10'h118 == io_rdAddr_0 ? lvtReg_280 : _GEN_4375; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4377 = 10'h119 == io_rdAddr_0 ? lvtReg_281 : _GEN_4376; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4378 = 10'h11a == io_rdAddr_0 ? lvtReg_282 : _GEN_4377; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4379 = 10'h11b == io_rdAddr_0 ? lvtReg_283 : _GEN_4378; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4380 = 10'h11c == io_rdAddr_0 ? lvtReg_284 : _GEN_4379; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4381 = 10'h11d == io_rdAddr_0 ? lvtReg_285 : _GEN_4380; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4382 = 10'h11e == io_rdAddr_0 ? lvtReg_286 : _GEN_4381; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4383 = 10'h11f == io_rdAddr_0 ? lvtReg_287 : _GEN_4382; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4384 = 10'h120 == io_rdAddr_0 ? lvtReg_288 : _GEN_4383; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4385 = 10'h121 == io_rdAddr_0 ? lvtReg_289 : _GEN_4384; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4386 = 10'h122 == io_rdAddr_0 ? lvtReg_290 : _GEN_4385; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4387 = 10'h123 == io_rdAddr_0 ? lvtReg_291 : _GEN_4386; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4388 = 10'h124 == io_rdAddr_0 ? lvtReg_292 : _GEN_4387; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4389 = 10'h125 == io_rdAddr_0 ? lvtReg_293 : _GEN_4388; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4390 = 10'h126 == io_rdAddr_0 ? lvtReg_294 : _GEN_4389; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4391 = 10'h127 == io_rdAddr_0 ? lvtReg_295 : _GEN_4390; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4392 = 10'h128 == io_rdAddr_0 ? lvtReg_296 : _GEN_4391; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4393 = 10'h129 == io_rdAddr_0 ? lvtReg_297 : _GEN_4392; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4394 = 10'h12a == io_rdAddr_0 ? lvtReg_298 : _GEN_4393; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4395 = 10'h12b == io_rdAddr_0 ? lvtReg_299 : _GEN_4394; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4396 = 10'h12c == io_rdAddr_0 ? lvtReg_300 : _GEN_4395; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4397 = 10'h12d == io_rdAddr_0 ? lvtReg_301 : _GEN_4396; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4398 = 10'h12e == io_rdAddr_0 ? lvtReg_302 : _GEN_4397; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4399 = 10'h12f == io_rdAddr_0 ? lvtReg_303 : _GEN_4398; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4400 = 10'h130 == io_rdAddr_0 ? lvtReg_304 : _GEN_4399; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4401 = 10'h131 == io_rdAddr_0 ? lvtReg_305 : _GEN_4400; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4402 = 10'h132 == io_rdAddr_0 ? lvtReg_306 : _GEN_4401; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4403 = 10'h133 == io_rdAddr_0 ? lvtReg_307 : _GEN_4402; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4404 = 10'h134 == io_rdAddr_0 ? lvtReg_308 : _GEN_4403; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4405 = 10'h135 == io_rdAddr_0 ? lvtReg_309 : _GEN_4404; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4406 = 10'h136 == io_rdAddr_0 ? lvtReg_310 : _GEN_4405; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4407 = 10'h137 == io_rdAddr_0 ? lvtReg_311 : _GEN_4406; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4408 = 10'h138 == io_rdAddr_0 ? lvtReg_312 : _GEN_4407; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4409 = 10'h139 == io_rdAddr_0 ? lvtReg_313 : _GEN_4408; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4410 = 10'h13a == io_rdAddr_0 ? lvtReg_314 : _GEN_4409; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4411 = 10'h13b == io_rdAddr_0 ? lvtReg_315 : _GEN_4410; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4412 = 10'h13c == io_rdAddr_0 ? lvtReg_316 : _GEN_4411; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4413 = 10'h13d == io_rdAddr_0 ? lvtReg_317 : _GEN_4412; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4414 = 10'h13e == io_rdAddr_0 ? lvtReg_318 : _GEN_4413; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4415 = 10'h13f == io_rdAddr_0 ? lvtReg_319 : _GEN_4414; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4416 = 10'h140 == io_rdAddr_0 ? lvtReg_320 : _GEN_4415; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4417 = 10'h141 == io_rdAddr_0 ? lvtReg_321 : _GEN_4416; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4418 = 10'h142 == io_rdAddr_0 ? lvtReg_322 : _GEN_4417; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4419 = 10'h143 == io_rdAddr_0 ? lvtReg_323 : _GEN_4418; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4420 = 10'h144 == io_rdAddr_0 ? lvtReg_324 : _GEN_4419; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4421 = 10'h145 == io_rdAddr_0 ? lvtReg_325 : _GEN_4420; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4422 = 10'h146 == io_rdAddr_0 ? lvtReg_326 : _GEN_4421; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4423 = 10'h147 == io_rdAddr_0 ? lvtReg_327 : _GEN_4422; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4424 = 10'h148 == io_rdAddr_0 ? lvtReg_328 : _GEN_4423; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4425 = 10'h149 == io_rdAddr_0 ? lvtReg_329 : _GEN_4424; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4426 = 10'h14a == io_rdAddr_0 ? lvtReg_330 : _GEN_4425; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4427 = 10'h14b == io_rdAddr_0 ? lvtReg_331 : _GEN_4426; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4428 = 10'h14c == io_rdAddr_0 ? lvtReg_332 : _GEN_4427; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4429 = 10'h14d == io_rdAddr_0 ? lvtReg_333 : _GEN_4428; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4430 = 10'h14e == io_rdAddr_0 ? lvtReg_334 : _GEN_4429; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4431 = 10'h14f == io_rdAddr_0 ? lvtReg_335 : _GEN_4430; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4432 = 10'h150 == io_rdAddr_0 ? lvtReg_336 : _GEN_4431; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4433 = 10'h151 == io_rdAddr_0 ? lvtReg_337 : _GEN_4432; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4434 = 10'h152 == io_rdAddr_0 ? lvtReg_338 : _GEN_4433; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4435 = 10'h153 == io_rdAddr_0 ? lvtReg_339 : _GEN_4434; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4436 = 10'h154 == io_rdAddr_0 ? lvtReg_340 : _GEN_4435; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4437 = 10'h155 == io_rdAddr_0 ? lvtReg_341 : _GEN_4436; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4438 = 10'h156 == io_rdAddr_0 ? lvtReg_342 : _GEN_4437; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4439 = 10'h157 == io_rdAddr_0 ? lvtReg_343 : _GEN_4438; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4440 = 10'h158 == io_rdAddr_0 ? lvtReg_344 : _GEN_4439; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4441 = 10'h159 == io_rdAddr_0 ? lvtReg_345 : _GEN_4440; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4442 = 10'h15a == io_rdAddr_0 ? lvtReg_346 : _GEN_4441; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4443 = 10'h15b == io_rdAddr_0 ? lvtReg_347 : _GEN_4442; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4444 = 10'h15c == io_rdAddr_0 ? lvtReg_348 : _GEN_4443; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4445 = 10'h15d == io_rdAddr_0 ? lvtReg_349 : _GEN_4444; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4446 = 10'h15e == io_rdAddr_0 ? lvtReg_350 : _GEN_4445; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4447 = 10'h15f == io_rdAddr_0 ? lvtReg_351 : _GEN_4446; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4448 = 10'h160 == io_rdAddr_0 ? lvtReg_352 : _GEN_4447; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4449 = 10'h161 == io_rdAddr_0 ? lvtReg_353 : _GEN_4448; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4450 = 10'h162 == io_rdAddr_0 ? lvtReg_354 : _GEN_4449; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4451 = 10'h163 == io_rdAddr_0 ? lvtReg_355 : _GEN_4450; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4452 = 10'h164 == io_rdAddr_0 ? lvtReg_356 : _GEN_4451; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4453 = 10'h165 == io_rdAddr_0 ? lvtReg_357 : _GEN_4452; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4454 = 10'h166 == io_rdAddr_0 ? lvtReg_358 : _GEN_4453; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4455 = 10'h167 == io_rdAddr_0 ? lvtReg_359 : _GEN_4454; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4456 = 10'h168 == io_rdAddr_0 ? lvtReg_360 : _GEN_4455; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4457 = 10'h169 == io_rdAddr_0 ? lvtReg_361 : _GEN_4456; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4458 = 10'h16a == io_rdAddr_0 ? lvtReg_362 : _GEN_4457; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4459 = 10'h16b == io_rdAddr_0 ? lvtReg_363 : _GEN_4458; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4460 = 10'h16c == io_rdAddr_0 ? lvtReg_364 : _GEN_4459; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4461 = 10'h16d == io_rdAddr_0 ? lvtReg_365 : _GEN_4460; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4462 = 10'h16e == io_rdAddr_0 ? lvtReg_366 : _GEN_4461; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4463 = 10'h16f == io_rdAddr_0 ? lvtReg_367 : _GEN_4462; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4464 = 10'h170 == io_rdAddr_0 ? lvtReg_368 : _GEN_4463; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4465 = 10'h171 == io_rdAddr_0 ? lvtReg_369 : _GEN_4464; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4466 = 10'h172 == io_rdAddr_0 ? lvtReg_370 : _GEN_4465; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4467 = 10'h173 == io_rdAddr_0 ? lvtReg_371 : _GEN_4466; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4468 = 10'h174 == io_rdAddr_0 ? lvtReg_372 : _GEN_4467; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4469 = 10'h175 == io_rdAddr_0 ? lvtReg_373 : _GEN_4468; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4470 = 10'h176 == io_rdAddr_0 ? lvtReg_374 : _GEN_4469; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4471 = 10'h177 == io_rdAddr_0 ? lvtReg_375 : _GEN_4470; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4472 = 10'h178 == io_rdAddr_0 ? lvtReg_376 : _GEN_4471; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4473 = 10'h179 == io_rdAddr_0 ? lvtReg_377 : _GEN_4472; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4474 = 10'h17a == io_rdAddr_0 ? lvtReg_378 : _GEN_4473; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4475 = 10'h17b == io_rdAddr_0 ? lvtReg_379 : _GEN_4474; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4476 = 10'h17c == io_rdAddr_0 ? lvtReg_380 : _GEN_4475; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4477 = 10'h17d == io_rdAddr_0 ? lvtReg_381 : _GEN_4476; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4478 = 10'h17e == io_rdAddr_0 ? lvtReg_382 : _GEN_4477; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4479 = 10'h17f == io_rdAddr_0 ? lvtReg_383 : _GEN_4478; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4480 = 10'h180 == io_rdAddr_0 ? lvtReg_384 : _GEN_4479; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4481 = 10'h181 == io_rdAddr_0 ? lvtReg_385 : _GEN_4480; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4482 = 10'h182 == io_rdAddr_0 ? lvtReg_386 : _GEN_4481; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4483 = 10'h183 == io_rdAddr_0 ? lvtReg_387 : _GEN_4482; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4484 = 10'h184 == io_rdAddr_0 ? lvtReg_388 : _GEN_4483; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4485 = 10'h185 == io_rdAddr_0 ? lvtReg_389 : _GEN_4484; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4486 = 10'h186 == io_rdAddr_0 ? lvtReg_390 : _GEN_4485; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4487 = 10'h187 == io_rdAddr_0 ? lvtReg_391 : _GEN_4486; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4488 = 10'h188 == io_rdAddr_0 ? lvtReg_392 : _GEN_4487; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4489 = 10'h189 == io_rdAddr_0 ? lvtReg_393 : _GEN_4488; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4490 = 10'h18a == io_rdAddr_0 ? lvtReg_394 : _GEN_4489; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4491 = 10'h18b == io_rdAddr_0 ? lvtReg_395 : _GEN_4490; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4492 = 10'h18c == io_rdAddr_0 ? lvtReg_396 : _GEN_4491; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4493 = 10'h18d == io_rdAddr_0 ? lvtReg_397 : _GEN_4492; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4494 = 10'h18e == io_rdAddr_0 ? lvtReg_398 : _GEN_4493; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4495 = 10'h18f == io_rdAddr_0 ? lvtReg_399 : _GEN_4494; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4496 = 10'h190 == io_rdAddr_0 ? lvtReg_400 : _GEN_4495; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4497 = 10'h191 == io_rdAddr_0 ? lvtReg_401 : _GEN_4496; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4498 = 10'h192 == io_rdAddr_0 ? lvtReg_402 : _GEN_4497; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4499 = 10'h193 == io_rdAddr_0 ? lvtReg_403 : _GEN_4498; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4500 = 10'h194 == io_rdAddr_0 ? lvtReg_404 : _GEN_4499; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4501 = 10'h195 == io_rdAddr_0 ? lvtReg_405 : _GEN_4500; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4502 = 10'h196 == io_rdAddr_0 ? lvtReg_406 : _GEN_4501; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4503 = 10'h197 == io_rdAddr_0 ? lvtReg_407 : _GEN_4502; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4504 = 10'h198 == io_rdAddr_0 ? lvtReg_408 : _GEN_4503; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4505 = 10'h199 == io_rdAddr_0 ? lvtReg_409 : _GEN_4504; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4506 = 10'h19a == io_rdAddr_0 ? lvtReg_410 : _GEN_4505; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4507 = 10'h19b == io_rdAddr_0 ? lvtReg_411 : _GEN_4506; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4508 = 10'h19c == io_rdAddr_0 ? lvtReg_412 : _GEN_4507; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4509 = 10'h19d == io_rdAddr_0 ? lvtReg_413 : _GEN_4508; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4510 = 10'h19e == io_rdAddr_0 ? lvtReg_414 : _GEN_4509; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4511 = 10'h19f == io_rdAddr_0 ? lvtReg_415 : _GEN_4510; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4512 = 10'h1a0 == io_rdAddr_0 ? lvtReg_416 : _GEN_4511; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4513 = 10'h1a1 == io_rdAddr_0 ? lvtReg_417 : _GEN_4512; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4514 = 10'h1a2 == io_rdAddr_0 ? lvtReg_418 : _GEN_4513; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4515 = 10'h1a3 == io_rdAddr_0 ? lvtReg_419 : _GEN_4514; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4516 = 10'h1a4 == io_rdAddr_0 ? lvtReg_420 : _GEN_4515; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4517 = 10'h1a5 == io_rdAddr_0 ? lvtReg_421 : _GEN_4516; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4518 = 10'h1a6 == io_rdAddr_0 ? lvtReg_422 : _GEN_4517; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4519 = 10'h1a7 == io_rdAddr_0 ? lvtReg_423 : _GEN_4518; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4520 = 10'h1a8 == io_rdAddr_0 ? lvtReg_424 : _GEN_4519; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4521 = 10'h1a9 == io_rdAddr_0 ? lvtReg_425 : _GEN_4520; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4522 = 10'h1aa == io_rdAddr_0 ? lvtReg_426 : _GEN_4521; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4523 = 10'h1ab == io_rdAddr_0 ? lvtReg_427 : _GEN_4522; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4524 = 10'h1ac == io_rdAddr_0 ? lvtReg_428 : _GEN_4523; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4525 = 10'h1ad == io_rdAddr_0 ? lvtReg_429 : _GEN_4524; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4526 = 10'h1ae == io_rdAddr_0 ? lvtReg_430 : _GEN_4525; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4527 = 10'h1af == io_rdAddr_0 ? lvtReg_431 : _GEN_4526; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4528 = 10'h1b0 == io_rdAddr_0 ? lvtReg_432 : _GEN_4527; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4529 = 10'h1b1 == io_rdAddr_0 ? lvtReg_433 : _GEN_4528; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4530 = 10'h1b2 == io_rdAddr_0 ? lvtReg_434 : _GEN_4529; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4531 = 10'h1b3 == io_rdAddr_0 ? lvtReg_435 : _GEN_4530; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4532 = 10'h1b4 == io_rdAddr_0 ? lvtReg_436 : _GEN_4531; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4533 = 10'h1b5 == io_rdAddr_0 ? lvtReg_437 : _GEN_4532; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4534 = 10'h1b6 == io_rdAddr_0 ? lvtReg_438 : _GEN_4533; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4535 = 10'h1b7 == io_rdAddr_0 ? lvtReg_439 : _GEN_4534; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4536 = 10'h1b8 == io_rdAddr_0 ? lvtReg_440 : _GEN_4535; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4537 = 10'h1b9 == io_rdAddr_0 ? lvtReg_441 : _GEN_4536; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4538 = 10'h1ba == io_rdAddr_0 ? lvtReg_442 : _GEN_4537; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4539 = 10'h1bb == io_rdAddr_0 ? lvtReg_443 : _GEN_4538; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4540 = 10'h1bc == io_rdAddr_0 ? lvtReg_444 : _GEN_4539; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4541 = 10'h1bd == io_rdAddr_0 ? lvtReg_445 : _GEN_4540; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4542 = 10'h1be == io_rdAddr_0 ? lvtReg_446 : _GEN_4541; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4543 = 10'h1bf == io_rdAddr_0 ? lvtReg_447 : _GEN_4542; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4544 = 10'h1c0 == io_rdAddr_0 ? lvtReg_448 : _GEN_4543; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4545 = 10'h1c1 == io_rdAddr_0 ? lvtReg_449 : _GEN_4544; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4546 = 10'h1c2 == io_rdAddr_0 ? lvtReg_450 : _GEN_4545; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4547 = 10'h1c3 == io_rdAddr_0 ? lvtReg_451 : _GEN_4546; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4548 = 10'h1c4 == io_rdAddr_0 ? lvtReg_452 : _GEN_4547; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4549 = 10'h1c5 == io_rdAddr_0 ? lvtReg_453 : _GEN_4548; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4550 = 10'h1c6 == io_rdAddr_0 ? lvtReg_454 : _GEN_4549; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4551 = 10'h1c7 == io_rdAddr_0 ? lvtReg_455 : _GEN_4550; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4552 = 10'h1c8 == io_rdAddr_0 ? lvtReg_456 : _GEN_4551; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4553 = 10'h1c9 == io_rdAddr_0 ? lvtReg_457 : _GEN_4552; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4554 = 10'h1ca == io_rdAddr_0 ? lvtReg_458 : _GEN_4553; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4555 = 10'h1cb == io_rdAddr_0 ? lvtReg_459 : _GEN_4554; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4556 = 10'h1cc == io_rdAddr_0 ? lvtReg_460 : _GEN_4555; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4557 = 10'h1cd == io_rdAddr_0 ? lvtReg_461 : _GEN_4556; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4558 = 10'h1ce == io_rdAddr_0 ? lvtReg_462 : _GEN_4557; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4559 = 10'h1cf == io_rdAddr_0 ? lvtReg_463 : _GEN_4558; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4560 = 10'h1d0 == io_rdAddr_0 ? lvtReg_464 : _GEN_4559; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4561 = 10'h1d1 == io_rdAddr_0 ? lvtReg_465 : _GEN_4560; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4562 = 10'h1d2 == io_rdAddr_0 ? lvtReg_466 : _GEN_4561; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4563 = 10'h1d3 == io_rdAddr_0 ? lvtReg_467 : _GEN_4562; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4564 = 10'h1d4 == io_rdAddr_0 ? lvtReg_468 : _GEN_4563; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4565 = 10'h1d5 == io_rdAddr_0 ? lvtReg_469 : _GEN_4564; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4566 = 10'h1d6 == io_rdAddr_0 ? lvtReg_470 : _GEN_4565; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4567 = 10'h1d7 == io_rdAddr_0 ? lvtReg_471 : _GEN_4566; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4568 = 10'h1d8 == io_rdAddr_0 ? lvtReg_472 : _GEN_4567; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4569 = 10'h1d9 == io_rdAddr_0 ? lvtReg_473 : _GEN_4568; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4570 = 10'h1da == io_rdAddr_0 ? lvtReg_474 : _GEN_4569; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4571 = 10'h1db == io_rdAddr_0 ? lvtReg_475 : _GEN_4570; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4572 = 10'h1dc == io_rdAddr_0 ? lvtReg_476 : _GEN_4571; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4573 = 10'h1dd == io_rdAddr_0 ? lvtReg_477 : _GEN_4572; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4574 = 10'h1de == io_rdAddr_0 ? lvtReg_478 : _GEN_4573; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4575 = 10'h1df == io_rdAddr_0 ? lvtReg_479 : _GEN_4574; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4576 = 10'h1e0 == io_rdAddr_0 ? lvtReg_480 : _GEN_4575; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4577 = 10'h1e1 == io_rdAddr_0 ? lvtReg_481 : _GEN_4576; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4578 = 10'h1e2 == io_rdAddr_0 ? lvtReg_482 : _GEN_4577; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4579 = 10'h1e3 == io_rdAddr_0 ? lvtReg_483 : _GEN_4578; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4580 = 10'h1e4 == io_rdAddr_0 ? lvtReg_484 : _GEN_4579; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4581 = 10'h1e5 == io_rdAddr_0 ? lvtReg_485 : _GEN_4580; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4582 = 10'h1e6 == io_rdAddr_0 ? lvtReg_486 : _GEN_4581; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4583 = 10'h1e7 == io_rdAddr_0 ? lvtReg_487 : _GEN_4582; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4584 = 10'h1e8 == io_rdAddr_0 ? lvtReg_488 : _GEN_4583; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4585 = 10'h1e9 == io_rdAddr_0 ? lvtReg_489 : _GEN_4584; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4586 = 10'h1ea == io_rdAddr_0 ? lvtReg_490 : _GEN_4585; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4587 = 10'h1eb == io_rdAddr_0 ? lvtReg_491 : _GEN_4586; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4588 = 10'h1ec == io_rdAddr_0 ? lvtReg_492 : _GEN_4587; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4589 = 10'h1ed == io_rdAddr_0 ? lvtReg_493 : _GEN_4588; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4590 = 10'h1ee == io_rdAddr_0 ? lvtReg_494 : _GEN_4589; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4591 = 10'h1ef == io_rdAddr_0 ? lvtReg_495 : _GEN_4590; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4592 = 10'h1f0 == io_rdAddr_0 ? lvtReg_496 : _GEN_4591; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4593 = 10'h1f1 == io_rdAddr_0 ? lvtReg_497 : _GEN_4592; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4594 = 10'h1f2 == io_rdAddr_0 ? lvtReg_498 : _GEN_4593; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4595 = 10'h1f3 == io_rdAddr_0 ? lvtReg_499 : _GEN_4594; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4596 = 10'h1f4 == io_rdAddr_0 ? lvtReg_500 : _GEN_4595; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4597 = 10'h1f5 == io_rdAddr_0 ? lvtReg_501 : _GEN_4596; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4598 = 10'h1f6 == io_rdAddr_0 ? lvtReg_502 : _GEN_4597; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4599 = 10'h1f7 == io_rdAddr_0 ? lvtReg_503 : _GEN_4598; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4600 = 10'h1f8 == io_rdAddr_0 ? lvtReg_504 : _GEN_4599; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4601 = 10'h1f9 == io_rdAddr_0 ? lvtReg_505 : _GEN_4600; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4602 = 10'h1fa == io_rdAddr_0 ? lvtReg_506 : _GEN_4601; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4603 = 10'h1fb == io_rdAddr_0 ? lvtReg_507 : _GEN_4602; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4604 = 10'h1fc == io_rdAddr_0 ? lvtReg_508 : _GEN_4603; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4605 = 10'h1fd == io_rdAddr_0 ? lvtReg_509 : _GEN_4604; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4606 = 10'h1fe == io_rdAddr_0 ? lvtReg_510 : _GEN_4605; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4607 = 10'h1ff == io_rdAddr_0 ? lvtReg_511 : _GEN_4606; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4608 = 10'h200 == io_rdAddr_0 ? lvtReg_512 : _GEN_4607; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4609 = 10'h201 == io_rdAddr_0 ? lvtReg_513 : _GEN_4608; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4610 = 10'h202 == io_rdAddr_0 ? lvtReg_514 : _GEN_4609; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4611 = 10'h203 == io_rdAddr_0 ? lvtReg_515 : _GEN_4610; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4612 = 10'h204 == io_rdAddr_0 ? lvtReg_516 : _GEN_4611; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4613 = 10'h205 == io_rdAddr_0 ? lvtReg_517 : _GEN_4612; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4614 = 10'h206 == io_rdAddr_0 ? lvtReg_518 : _GEN_4613; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4615 = 10'h207 == io_rdAddr_0 ? lvtReg_519 : _GEN_4614; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4616 = 10'h208 == io_rdAddr_0 ? lvtReg_520 : _GEN_4615; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4617 = 10'h209 == io_rdAddr_0 ? lvtReg_521 : _GEN_4616; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4618 = 10'h20a == io_rdAddr_0 ? lvtReg_522 : _GEN_4617; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4619 = 10'h20b == io_rdAddr_0 ? lvtReg_523 : _GEN_4618; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4620 = 10'h20c == io_rdAddr_0 ? lvtReg_524 : _GEN_4619; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4621 = 10'h20d == io_rdAddr_0 ? lvtReg_525 : _GEN_4620; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4622 = 10'h20e == io_rdAddr_0 ? lvtReg_526 : _GEN_4621; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4623 = 10'h20f == io_rdAddr_0 ? lvtReg_527 : _GEN_4622; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4624 = 10'h210 == io_rdAddr_0 ? lvtReg_528 : _GEN_4623; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4625 = 10'h211 == io_rdAddr_0 ? lvtReg_529 : _GEN_4624; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4626 = 10'h212 == io_rdAddr_0 ? lvtReg_530 : _GEN_4625; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4627 = 10'h213 == io_rdAddr_0 ? lvtReg_531 : _GEN_4626; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4628 = 10'h214 == io_rdAddr_0 ? lvtReg_532 : _GEN_4627; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4629 = 10'h215 == io_rdAddr_0 ? lvtReg_533 : _GEN_4628; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4630 = 10'h216 == io_rdAddr_0 ? lvtReg_534 : _GEN_4629; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4631 = 10'h217 == io_rdAddr_0 ? lvtReg_535 : _GEN_4630; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4632 = 10'h218 == io_rdAddr_0 ? lvtReg_536 : _GEN_4631; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4633 = 10'h219 == io_rdAddr_0 ? lvtReg_537 : _GEN_4632; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4634 = 10'h21a == io_rdAddr_0 ? lvtReg_538 : _GEN_4633; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4635 = 10'h21b == io_rdAddr_0 ? lvtReg_539 : _GEN_4634; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4636 = 10'h21c == io_rdAddr_0 ? lvtReg_540 : _GEN_4635; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4637 = 10'h21d == io_rdAddr_0 ? lvtReg_541 : _GEN_4636; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4638 = 10'h21e == io_rdAddr_0 ? lvtReg_542 : _GEN_4637; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4639 = 10'h21f == io_rdAddr_0 ? lvtReg_543 : _GEN_4638; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4640 = 10'h220 == io_rdAddr_0 ? lvtReg_544 : _GEN_4639; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4641 = 10'h221 == io_rdAddr_0 ? lvtReg_545 : _GEN_4640; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4642 = 10'h222 == io_rdAddr_0 ? lvtReg_546 : _GEN_4641; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4643 = 10'h223 == io_rdAddr_0 ? lvtReg_547 : _GEN_4642; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4644 = 10'h224 == io_rdAddr_0 ? lvtReg_548 : _GEN_4643; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4645 = 10'h225 == io_rdAddr_0 ? lvtReg_549 : _GEN_4644; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4646 = 10'h226 == io_rdAddr_0 ? lvtReg_550 : _GEN_4645; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4647 = 10'h227 == io_rdAddr_0 ? lvtReg_551 : _GEN_4646; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4648 = 10'h228 == io_rdAddr_0 ? lvtReg_552 : _GEN_4647; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4649 = 10'h229 == io_rdAddr_0 ? lvtReg_553 : _GEN_4648; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4650 = 10'h22a == io_rdAddr_0 ? lvtReg_554 : _GEN_4649; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4651 = 10'h22b == io_rdAddr_0 ? lvtReg_555 : _GEN_4650; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4652 = 10'h22c == io_rdAddr_0 ? lvtReg_556 : _GEN_4651; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4653 = 10'h22d == io_rdAddr_0 ? lvtReg_557 : _GEN_4652; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4654 = 10'h22e == io_rdAddr_0 ? lvtReg_558 : _GEN_4653; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4655 = 10'h22f == io_rdAddr_0 ? lvtReg_559 : _GEN_4654; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4656 = 10'h230 == io_rdAddr_0 ? lvtReg_560 : _GEN_4655; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4657 = 10'h231 == io_rdAddr_0 ? lvtReg_561 : _GEN_4656; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4658 = 10'h232 == io_rdAddr_0 ? lvtReg_562 : _GEN_4657; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4659 = 10'h233 == io_rdAddr_0 ? lvtReg_563 : _GEN_4658; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4660 = 10'h234 == io_rdAddr_0 ? lvtReg_564 : _GEN_4659; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4661 = 10'h235 == io_rdAddr_0 ? lvtReg_565 : _GEN_4660; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4662 = 10'h236 == io_rdAddr_0 ? lvtReg_566 : _GEN_4661; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4663 = 10'h237 == io_rdAddr_0 ? lvtReg_567 : _GEN_4662; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4664 = 10'h238 == io_rdAddr_0 ? lvtReg_568 : _GEN_4663; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4665 = 10'h239 == io_rdAddr_0 ? lvtReg_569 : _GEN_4664; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4666 = 10'h23a == io_rdAddr_0 ? lvtReg_570 : _GEN_4665; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4667 = 10'h23b == io_rdAddr_0 ? lvtReg_571 : _GEN_4666; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4668 = 10'h23c == io_rdAddr_0 ? lvtReg_572 : _GEN_4667; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4669 = 10'h23d == io_rdAddr_0 ? lvtReg_573 : _GEN_4668; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4670 = 10'h23e == io_rdAddr_0 ? lvtReg_574 : _GEN_4669; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4671 = 10'h23f == io_rdAddr_0 ? lvtReg_575 : _GEN_4670; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4672 = 10'h240 == io_rdAddr_0 ? lvtReg_576 : _GEN_4671; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4673 = 10'h241 == io_rdAddr_0 ? lvtReg_577 : _GEN_4672; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4674 = 10'h242 == io_rdAddr_0 ? lvtReg_578 : _GEN_4673; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4675 = 10'h243 == io_rdAddr_0 ? lvtReg_579 : _GEN_4674; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4676 = 10'h244 == io_rdAddr_0 ? lvtReg_580 : _GEN_4675; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4677 = 10'h245 == io_rdAddr_0 ? lvtReg_581 : _GEN_4676; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4678 = 10'h246 == io_rdAddr_0 ? lvtReg_582 : _GEN_4677; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4679 = 10'h247 == io_rdAddr_0 ? lvtReg_583 : _GEN_4678; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4680 = 10'h248 == io_rdAddr_0 ? lvtReg_584 : _GEN_4679; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4681 = 10'h249 == io_rdAddr_0 ? lvtReg_585 : _GEN_4680; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4682 = 10'h24a == io_rdAddr_0 ? lvtReg_586 : _GEN_4681; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4683 = 10'h24b == io_rdAddr_0 ? lvtReg_587 : _GEN_4682; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4684 = 10'h24c == io_rdAddr_0 ? lvtReg_588 : _GEN_4683; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4685 = 10'h24d == io_rdAddr_0 ? lvtReg_589 : _GEN_4684; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4686 = 10'h24e == io_rdAddr_0 ? lvtReg_590 : _GEN_4685; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4687 = 10'h24f == io_rdAddr_0 ? lvtReg_591 : _GEN_4686; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4688 = 10'h250 == io_rdAddr_0 ? lvtReg_592 : _GEN_4687; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4689 = 10'h251 == io_rdAddr_0 ? lvtReg_593 : _GEN_4688; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4690 = 10'h252 == io_rdAddr_0 ? lvtReg_594 : _GEN_4689; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4691 = 10'h253 == io_rdAddr_0 ? lvtReg_595 : _GEN_4690; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4692 = 10'h254 == io_rdAddr_0 ? lvtReg_596 : _GEN_4691; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4693 = 10'h255 == io_rdAddr_0 ? lvtReg_597 : _GEN_4692; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4694 = 10'h256 == io_rdAddr_0 ? lvtReg_598 : _GEN_4693; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4695 = 10'h257 == io_rdAddr_0 ? lvtReg_599 : _GEN_4694; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4696 = 10'h258 == io_rdAddr_0 ? lvtReg_600 : _GEN_4695; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4697 = 10'h259 == io_rdAddr_0 ? lvtReg_601 : _GEN_4696; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4698 = 10'h25a == io_rdAddr_0 ? lvtReg_602 : _GEN_4697; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4699 = 10'h25b == io_rdAddr_0 ? lvtReg_603 : _GEN_4698; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4700 = 10'h25c == io_rdAddr_0 ? lvtReg_604 : _GEN_4699; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4701 = 10'h25d == io_rdAddr_0 ? lvtReg_605 : _GEN_4700; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4702 = 10'h25e == io_rdAddr_0 ? lvtReg_606 : _GEN_4701; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4703 = 10'h25f == io_rdAddr_0 ? lvtReg_607 : _GEN_4702; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4704 = 10'h260 == io_rdAddr_0 ? lvtReg_608 : _GEN_4703; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4705 = 10'h261 == io_rdAddr_0 ? lvtReg_609 : _GEN_4704; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4706 = 10'h262 == io_rdAddr_0 ? lvtReg_610 : _GEN_4705; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4707 = 10'h263 == io_rdAddr_0 ? lvtReg_611 : _GEN_4706; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4708 = 10'h264 == io_rdAddr_0 ? lvtReg_612 : _GEN_4707; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4709 = 10'h265 == io_rdAddr_0 ? lvtReg_613 : _GEN_4708; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4710 = 10'h266 == io_rdAddr_0 ? lvtReg_614 : _GEN_4709; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4711 = 10'h267 == io_rdAddr_0 ? lvtReg_615 : _GEN_4710; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4712 = 10'h268 == io_rdAddr_0 ? lvtReg_616 : _GEN_4711; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4713 = 10'h269 == io_rdAddr_0 ? lvtReg_617 : _GEN_4712; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4714 = 10'h26a == io_rdAddr_0 ? lvtReg_618 : _GEN_4713; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4715 = 10'h26b == io_rdAddr_0 ? lvtReg_619 : _GEN_4714; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4716 = 10'h26c == io_rdAddr_0 ? lvtReg_620 : _GEN_4715; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4717 = 10'h26d == io_rdAddr_0 ? lvtReg_621 : _GEN_4716; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4718 = 10'h26e == io_rdAddr_0 ? lvtReg_622 : _GEN_4717; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4719 = 10'h26f == io_rdAddr_0 ? lvtReg_623 : _GEN_4718; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4720 = 10'h270 == io_rdAddr_0 ? lvtReg_624 : _GEN_4719; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4721 = 10'h271 == io_rdAddr_0 ? lvtReg_625 : _GEN_4720; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4722 = 10'h272 == io_rdAddr_0 ? lvtReg_626 : _GEN_4721; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4723 = 10'h273 == io_rdAddr_0 ? lvtReg_627 : _GEN_4722; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4724 = 10'h274 == io_rdAddr_0 ? lvtReg_628 : _GEN_4723; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4725 = 10'h275 == io_rdAddr_0 ? lvtReg_629 : _GEN_4724; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4726 = 10'h276 == io_rdAddr_0 ? lvtReg_630 : _GEN_4725; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4727 = 10'h277 == io_rdAddr_0 ? lvtReg_631 : _GEN_4726; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4728 = 10'h278 == io_rdAddr_0 ? lvtReg_632 : _GEN_4727; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4729 = 10'h279 == io_rdAddr_0 ? lvtReg_633 : _GEN_4728; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4730 = 10'h27a == io_rdAddr_0 ? lvtReg_634 : _GEN_4729; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4731 = 10'h27b == io_rdAddr_0 ? lvtReg_635 : _GEN_4730; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4732 = 10'h27c == io_rdAddr_0 ? lvtReg_636 : _GEN_4731; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4733 = 10'h27d == io_rdAddr_0 ? lvtReg_637 : _GEN_4732; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4734 = 10'h27e == io_rdAddr_0 ? lvtReg_638 : _GEN_4733; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4735 = 10'h27f == io_rdAddr_0 ? lvtReg_639 : _GEN_4734; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4736 = 10'h280 == io_rdAddr_0 ? lvtReg_640 : _GEN_4735; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4737 = 10'h281 == io_rdAddr_0 ? lvtReg_641 : _GEN_4736; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4738 = 10'h282 == io_rdAddr_0 ? lvtReg_642 : _GEN_4737; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4739 = 10'h283 == io_rdAddr_0 ? lvtReg_643 : _GEN_4738; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4740 = 10'h284 == io_rdAddr_0 ? lvtReg_644 : _GEN_4739; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4741 = 10'h285 == io_rdAddr_0 ? lvtReg_645 : _GEN_4740; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4742 = 10'h286 == io_rdAddr_0 ? lvtReg_646 : _GEN_4741; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4743 = 10'h287 == io_rdAddr_0 ? lvtReg_647 : _GEN_4742; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4744 = 10'h288 == io_rdAddr_0 ? lvtReg_648 : _GEN_4743; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4745 = 10'h289 == io_rdAddr_0 ? lvtReg_649 : _GEN_4744; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4746 = 10'h28a == io_rdAddr_0 ? lvtReg_650 : _GEN_4745; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4747 = 10'h28b == io_rdAddr_0 ? lvtReg_651 : _GEN_4746; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4748 = 10'h28c == io_rdAddr_0 ? lvtReg_652 : _GEN_4747; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4749 = 10'h28d == io_rdAddr_0 ? lvtReg_653 : _GEN_4748; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4750 = 10'h28e == io_rdAddr_0 ? lvtReg_654 : _GEN_4749; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4751 = 10'h28f == io_rdAddr_0 ? lvtReg_655 : _GEN_4750; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4752 = 10'h290 == io_rdAddr_0 ? lvtReg_656 : _GEN_4751; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4753 = 10'h291 == io_rdAddr_0 ? lvtReg_657 : _GEN_4752; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4754 = 10'h292 == io_rdAddr_0 ? lvtReg_658 : _GEN_4753; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4755 = 10'h293 == io_rdAddr_0 ? lvtReg_659 : _GEN_4754; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4756 = 10'h294 == io_rdAddr_0 ? lvtReg_660 : _GEN_4755; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4757 = 10'h295 == io_rdAddr_0 ? lvtReg_661 : _GEN_4756; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4758 = 10'h296 == io_rdAddr_0 ? lvtReg_662 : _GEN_4757; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4759 = 10'h297 == io_rdAddr_0 ? lvtReg_663 : _GEN_4758; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4760 = 10'h298 == io_rdAddr_0 ? lvtReg_664 : _GEN_4759; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4761 = 10'h299 == io_rdAddr_0 ? lvtReg_665 : _GEN_4760; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4762 = 10'h29a == io_rdAddr_0 ? lvtReg_666 : _GEN_4761; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4763 = 10'h29b == io_rdAddr_0 ? lvtReg_667 : _GEN_4762; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4764 = 10'h29c == io_rdAddr_0 ? lvtReg_668 : _GEN_4763; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4765 = 10'h29d == io_rdAddr_0 ? lvtReg_669 : _GEN_4764; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4766 = 10'h29e == io_rdAddr_0 ? lvtReg_670 : _GEN_4765; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4767 = 10'h29f == io_rdAddr_0 ? lvtReg_671 : _GEN_4766; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4768 = 10'h2a0 == io_rdAddr_0 ? lvtReg_672 : _GEN_4767; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4769 = 10'h2a1 == io_rdAddr_0 ? lvtReg_673 : _GEN_4768; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4770 = 10'h2a2 == io_rdAddr_0 ? lvtReg_674 : _GEN_4769; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4771 = 10'h2a3 == io_rdAddr_0 ? lvtReg_675 : _GEN_4770; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4772 = 10'h2a4 == io_rdAddr_0 ? lvtReg_676 : _GEN_4771; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4773 = 10'h2a5 == io_rdAddr_0 ? lvtReg_677 : _GEN_4772; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4774 = 10'h2a6 == io_rdAddr_0 ? lvtReg_678 : _GEN_4773; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4775 = 10'h2a7 == io_rdAddr_0 ? lvtReg_679 : _GEN_4774; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4776 = 10'h2a8 == io_rdAddr_0 ? lvtReg_680 : _GEN_4775; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4777 = 10'h2a9 == io_rdAddr_0 ? lvtReg_681 : _GEN_4776; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4778 = 10'h2aa == io_rdAddr_0 ? lvtReg_682 : _GEN_4777; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4779 = 10'h2ab == io_rdAddr_0 ? lvtReg_683 : _GEN_4778; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4780 = 10'h2ac == io_rdAddr_0 ? lvtReg_684 : _GEN_4779; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4781 = 10'h2ad == io_rdAddr_0 ? lvtReg_685 : _GEN_4780; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4782 = 10'h2ae == io_rdAddr_0 ? lvtReg_686 : _GEN_4781; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4783 = 10'h2af == io_rdAddr_0 ? lvtReg_687 : _GEN_4782; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4784 = 10'h2b0 == io_rdAddr_0 ? lvtReg_688 : _GEN_4783; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4785 = 10'h2b1 == io_rdAddr_0 ? lvtReg_689 : _GEN_4784; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4786 = 10'h2b2 == io_rdAddr_0 ? lvtReg_690 : _GEN_4785; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4787 = 10'h2b3 == io_rdAddr_0 ? lvtReg_691 : _GEN_4786; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4788 = 10'h2b4 == io_rdAddr_0 ? lvtReg_692 : _GEN_4787; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4789 = 10'h2b5 == io_rdAddr_0 ? lvtReg_693 : _GEN_4788; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4790 = 10'h2b6 == io_rdAddr_0 ? lvtReg_694 : _GEN_4789; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4791 = 10'h2b7 == io_rdAddr_0 ? lvtReg_695 : _GEN_4790; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4792 = 10'h2b8 == io_rdAddr_0 ? lvtReg_696 : _GEN_4791; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4793 = 10'h2b9 == io_rdAddr_0 ? lvtReg_697 : _GEN_4792; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4794 = 10'h2ba == io_rdAddr_0 ? lvtReg_698 : _GEN_4793; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4795 = 10'h2bb == io_rdAddr_0 ? lvtReg_699 : _GEN_4794; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4796 = 10'h2bc == io_rdAddr_0 ? lvtReg_700 : _GEN_4795; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4797 = 10'h2bd == io_rdAddr_0 ? lvtReg_701 : _GEN_4796; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4798 = 10'h2be == io_rdAddr_0 ? lvtReg_702 : _GEN_4797; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4799 = 10'h2bf == io_rdAddr_0 ? lvtReg_703 : _GEN_4798; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4800 = 10'h2c0 == io_rdAddr_0 ? lvtReg_704 : _GEN_4799; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4801 = 10'h2c1 == io_rdAddr_0 ? lvtReg_705 : _GEN_4800; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4802 = 10'h2c2 == io_rdAddr_0 ? lvtReg_706 : _GEN_4801; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4803 = 10'h2c3 == io_rdAddr_0 ? lvtReg_707 : _GEN_4802; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4804 = 10'h2c4 == io_rdAddr_0 ? lvtReg_708 : _GEN_4803; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4805 = 10'h2c5 == io_rdAddr_0 ? lvtReg_709 : _GEN_4804; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4806 = 10'h2c6 == io_rdAddr_0 ? lvtReg_710 : _GEN_4805; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4807 = 10'h2c7 == io_rdAddr_0 ? lvtReg_711 : _GEN_4806; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4808 = 10'h2c8 == io_rdAddr_0 ? lvtReg_712 : _GEN_4807; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4809 = 10'h2c9 == io_rdAddr_0 ? lvtReg_713 : _GEN_4808; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4810 = 10'h2ca == io_rdAddr_0 ? lvtReg_714 : _GEN_4809; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4811 = 10'h2cb == io_rdAddr_0 ? lvtReg_715 : _GEN_4810; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4812 = 10'h2cc == io_rdAddr_0 ? lvtReg_716 : _GEN_4811; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4813 = 10'h2cd == io_rdAddr_0 ? lvtReg_717 : _GEN_4812; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4814 = 10'h2ce == io_rdAddr_0 ? lvtReg_718 : _GEN_4813; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4815 = 10'h2cf == io_rdAddr_0 ? lvtReg_719 : _GEN_4814; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4816 = 10'h2d0 == io_rdAddr_0 ? lvtReg_720 : _GEN_4815; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4817 = 10'h2d1 == io_rdAddr_0 ? lvtReg_721 : _GEN_4816; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4818 = 10'h2d2 == io_rdAddr_0 ? lvtReg_722 : _GEN_4817; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4819 = 10'h2d3 == io_rdAddr_0 ? lvtReg_723 : _GEN_4818; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4820 = 10'h2d4 == io_rdAddr_0 ? lvtReg_724 : _GEN_4819; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4821 = 10'h2d5 == io_rdAddr_0 ? lvtReg_725 : _GEN_4820; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4822 = 10'h2d6 == io_rdAddr_0 ? lvtReg_726 : _GEN_4821; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4823 = 10'h2d7 == io_rdAddr_0 ? lvtReg_727 : _GEN_4822; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4824 = 10'h2d8 == io_rdAddr_0 ? lvtReg_728 : _GEN_4823; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4825 = 10'h2d9 == io_rdAddr_0 ? lvtReg_729 : _GEN_4824; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4826 = 10'h2da == io_rdAddr_0 ? lvtReg_730 : _GEN_4825; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4827 = 10'h2db == io_rdAddr_0 ? lvtReg_731 : _GEN_4826; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4828 = 10'h2dc == io_rdAddr_0 ? lvtReg_732 : _GEN_4827; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4829 = 10'h2dd == io_rdAddr_0 ? lvtReg_733 : _GEN_4828; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4830 = 10'h2de == io_rdAddr_0 ? lvtReg_734 : _GEN_4829; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4831 = 10'h2df == io_rdAddr_0 ? lvtReg_735 : _GEN_4830; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4832 = 10'h2e0 == io_rdAddr_0 ? lvtReg_736 : _GEN_4831; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4833 = 10'h2e1 == io_rdAddr_0 ? lvtReg_737 : _GEN_4832; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4834 = 10'h2e2 == io_rdAddr_0 ? lvtReg_738 : _GEN_4833; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4835 = 10'h2e3 == io_rdAddr_0 ? lvtReg_739 : _GEN_4834; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4836 = 10'h2e4 == io_rdAddr_0 ? lvtReg_740 : _GEN_4835; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4837 = 10'h2e5 == io_rdAddr_0 ? lvtReg_741 : _GEN_4836; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4838 = 10'h2e6 == io_rdAddr_0 ? lvtReg_742 : _GEN_4837; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4839 = 10'h2e7 == io_rdAddr_0 ? lvtReg_743 : _GEN_4838; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4840 = 10'h2e8 == io_rdAddr_0 ? lvtReg_744 : _GEN_4839; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4841 = 10'h2e9 == io_rdAddr_0 ? lvtReg_745 : _GEN_4840; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4842 = 10'h2ea == io_rdAddr_0 ? lvtReg_746 : _GEN_4841; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4843 = 10'h2eb == io_rdAddr_0 ? lvtReg_747 : _GEN_4842; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4844 = 10'h2ec == io_rdAddr_0 ? lvtReg_748 : _GEN_4843; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4845 = 10'h2ed == io_rdAddr_0 ? lvtReg_749 : _GEN_4844; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4846 = 10'h2ee == io_rdAddr_0 ? lvtReg_750 : _GEN_4845; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4847 = 10'h2ef == io_rdAddr_0 ? lvtReg_751 : _GEN_4846; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4848 = 10'h2f0 == io_rdAddr_0 ? lvtReg_752 : _GEN_4847; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4849 = 10'h2f1 == io_rdAddr_0 ? lvtReg_753 : _GEN_4848; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4850 = 10'h2f2 == io_rdAddr_0 ? lvtReg_754 : _GEN_4849; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4851 = 10'h2f3 == io_rdAddr_0 ? lvtReg_755 : _GEN_4850; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4852 = 10'h2f4 == io_rdAddr_0 ? lvtReg_756 : _GEN_4851; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4853 = 10'h2f5 == io_rdAddr_0 ? lvtReg_757 : _GEN_4852; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4854 = 10'h2f6 == io_rdAddr_0 ? lvtReg_758 : _GEN_4853; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4855 = 10'h2f7 == io_rdAddr_0 ? lvtReg_759 : _GEN_4854; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4856 = 10'h2f8 == io_rdAddr_0 ? lvtReg_760 : _GEN_4855; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4857 = 10'h2f9 == io_rdAddr_0 ? lvtReg_761 : _GEN_4856; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4858 = 10'h2fa == io_rdAddr_0 ? lvtReg_762 : _GEN_4857; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4859 = 10'h2fb == io_rdAddr_0 ? lvtReg_763 : _GEN_4858; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4860 = 10'h2fc == io_rdAddr_0 ? lvtReg_764 : _GEN_4859; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4861 = 10'h2fd == io_rdAddr_0 ? lvtReg_765 : _GEN_4860; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4862 = 10'h2fe == io_rdAddr_0 ? lvtReg_766 : _GEN_4861; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4863 = 10'h2ff == io_rdAddr_0 ? lvtReg_767 : _GEN_4862; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4864 = 10'h300 == io_rdAddr_0 ? lvtReg_768 : _GEN_4863; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4865 = 10'h301 == io_rdAddr_0 ? lvtReg_769 : _GEN_4864; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4866 = 10'h302 == io_rdAddr_0 ? lvtReg_770 : _GEN_4865; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4867 = 10'h303 == io_rdAddr_0 ? lvtReg_771 : _GEN_4866; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4868 = 10'h304 == io_rdAddr_0 ? lvtReg_772 : _GEN_4867; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4869 = 10'h305 == io_rdAddr_0 ? lvtReg_773 : _GEN_4868; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4870 = 10'h306 == io_rdAddr_0 ? lvtReg_774 : _GEN_4869; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4871 = 10'h307 == io_rdAddr_0 ? lvtReg_775 : _GEN_4870; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4872 = 10'h308 == io_rdAddr_0 ? lvtReg_776 : _GEN_4871; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4873 = 10'h309 == io_rdAddr_0 ? lvtReg_777 : _GEN_4872; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4874 = 10'h30a == io_rdAddr_0 ? lvtReg_778 : _GEN_4873; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4875 = 10'h30b == io_rdAddr_0 ? lvtReg_779 : _GEN_4874; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4876 = 10'h30c == io_rdAddr_0 ? lvtReg_780 : _GEN_4875; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4877 = 10'h30d == io_rdAddr_0 ? lvtReg_781 : _GEN_4876; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4878 = 10'h30e == io_rdAddr_0 ? lvtReg_782 : _GEN_4877; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4879 = 10'h30f == io_rdAddr_0 ? lvtReg_783 : _GEN_4878; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4880 = 10'h310 == io_rdAddr_0 ? lvtReg_784 : _GEN_4879; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4881 = 10'h311 == io_rdAddr_0 ? lvtReg_785 : _GEN_4880; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4882 = 10'h312 == io_rdAddr_0 ? lvtReg_786 : _GEN_4881; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4883 = 10'h313 == io_rdAddr_0 ? lvtReg_787 : _GEN_4882; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4884 = 10'h314 == io_rdAddr_0 ? lvtReg_788 : _GEN_4883; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4885 = 10'h315 == io_rdAddr_0 ? lvtReg_789 : _GEN_4884; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4886 = 10'h316 == io_rdAddr_0 ? lvtReg_790 : _GEN_4885; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4887 = 10'h317 == io_rdAddr_0 ? lvtReg_791 : _GEN_4886; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4888 = 10'h318 == io_rdAddr_0 ? lvtReg_792 : _GEN_4887; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4889 = 10'h319 == io_rdAddr_0 ? lvtReg_793 : _GEN_4888; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4890 = 10'h31a == io_rdAddr_0 ? lvtReg_794 : _GEN_4889; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4891 = 10'h31b == io_rdAddr_0 ? lvtReg_795 : _GEN_4890; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4892 = 10'h31c == io_rdAddr_0 ? lvtReg_796 : _GEN_4891; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4893 = 10'h31d == io_rdAddr_0 ? lvtReg_797 : _GEN_4892; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4894 = 10'h31e == io_rdAddr_0 ? lvtReg_798 : _GEN_4893; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4895 = 10'h31f == io_rdAddr_0 ? lvtReg_799 : _GEN_4894; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4896 = 10'h320 == io_rdAddr_0 ? lvtReg_800 : _GEN_4895; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4897 = 10'h321 == io_rdAddr_0 ? lvtReg_801 : _GEN_4896; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4898 = 10'h322 == io_rdAddr_0 ? lvtReg_802 : _GEN_4897; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4899 = 10'h323 == io_rdAddr_0 ? lvtReg_803 : _GEN_4898; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4900 = 10'h324 == io_rdAddr_0 ? lvtReg_804 : _GEN_4899; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4901 = 10'h325 == io_rdAddr_0 ? lvtReg_805 : _GEN_4900; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4902 = 10'h326 == io_rdAddr_0 ? lvtReg_806 : _GEN_4901; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4903 = 10'h327 == io_rdAddr_0 ? lvtReg_807 : _GEN_4902; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4904 = 10'h328 == io_rdAddr_0 ? lvtReg_808 : _GEN_4903; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4905 = 10'h329 == io_rdAddr_0 ? lvtReg_809 : _GEN_4904; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4906 = 10'h32a == io_rdAddr_0 ? lvtReg_810 : _GEN_4905; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4907 = 10'h32b == io_rdAddr_0 ? lvtReg_811 : _GEN_4906; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4908 = 10'h32c == io_rdAddr_0 ? lvtReg_812 : _GEN_4907; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4909 = 10'h32d == io_rdAddr_0 ? lvtReg_813 : _GEN_4908; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4910 = 10'h32e == io_rdAddr_0 ? lvtReg_814 : _GEN_4909; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4911 = 10'h32f == io_rdAddr_0 ? lvtReg_815 : _GEN_4910; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4912 = 10'h330 == io_rdAddr_0 ? lvtReg_816 : _GEN_4911; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4913 = 10'h331 == io_rdAddr_0 ? lvtReg_817 : _GEN_4912; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4914 = 10'h332 == io_rdAddr_0 ? lvtReg_818 : _GEN_4913; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4915 = 10'h333 == io_rdAddr_0 ? lvtReg_819 : _GEN_4914; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4916 = 10'h334 == io_rdAddr_0 ? lvtReg_820 : _GEN_4915; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4917 = 10'h335 == io_rdAddr_0 ? lvtReg_821 : _GEN_4916; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4918 = 10'h336 == io_rdAddr_0 ? lvtReg_822 : _GEN_4917; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4919 = 10'h337 == io_rdAddr_0 ? lvtReg_823 : _GEN_4918; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4920 = 10'h338 == io_rdAddr_0 ? lvtReg_824 : _GEN_4919; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4921 = 10'h339 == io_rdAddr_0 ? lvtReg_825 : _GEN_4920; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4922 = 10'h33a == io_rdAddr_0 ? lvtReg_826 : _GEN_4921; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4923 = 10'h33b == io_rdAddr_0 ? lvtReg_827 : _GEN_4922; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4924 = 10'h33c == io_rdAddr_0 ? lvtReg_828 : _GEN_4923; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4925 = 10'h33d == io_rdAddr_0 ? lvtReg_829 : _GEN_4924; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4926 = 10'h33e == io_rdAddr_0 ? lvtReg_830 : _GEN_4925; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4927 = 10'h33f == io_rdAddr_0 ? lvtReg_831 : _GEN_4926; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4928 = 10'h340 == io_rdAddr_0 ? lvtReg_832 : _GEN_4927; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4929 = 10'h341 == io_rdAddr_0 ? lvtReg_833 : _GEN_4928; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4930 = 10'h342 == io_rdAddr_0 ? lvtReg_834 : _GEN_4929; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4931 = 10'h343 == io_rdAddr_0 ? lvtReg_835 : _GEN_4930; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4932 = 10'h344 == io_rdAddr_0 ? lvtReg_836 : _GEN_4931; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4933 = 10'h345 == io_rdAddr_0 ? lvtReg_837 : _GEN_4932; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4934 = 10'h346 == io_rdAddr_0 ? lvtReg_838 : _GEN_4933; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4935 = 10'h347 == io_rdAddr_0 ? lvtReg_839 : _GEN_4934; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4936 = 10'h348 == io_rdAddr_0 ? lvtReg_840 : _GEN_4935; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4937 = 10'h349 == io_rdAddr_0 ? lvtReg_841 : _GEN_4936; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4938 = 10'h34a == io_rdAddr_0 ? lvtReg_842 : _GEN_4937; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4939 = 10'h34b == io_rdAddr_0 ? lvtReg_843 : _GEN_4938; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4940 = 10'h34c == io_rdAddr_0 ? lvtReg_844 : _GEN_4939; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4941 = 10'h34d == io_rdAddr_0 ? lvtReg_845 : _GEN_4940; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4942 = 10'h34e == io_rdAddr_0 ? lvtReg_846 : _GEN_4941; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4943 = 10'h34f == io_rdAddr_0 ? lvtReg_847 : _GEN_4942; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4944 = 10'h350 == io_rdAddr_0 ? lvtReg_848 : _GEN_4943; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4945 = 10'h351 == io_rdAddr_0 ? lvtReg_849 : _GEN_4944; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4946 = 10'h352 == io_rdAddr_0 ? lvtReg_850 : _GEN_4945; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4947 = 10'h353 == io_rdAddr_0 ? lvtReg_851 : _GEN_4946; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4948 = 10'h354 == io_rdAddr_0 ? lvtReg_852 : _GEN_4947; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4949 = 10'h355 == io_rdAddr_0 ? lvtReg_853 : _GEN_4948; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4950 = 10'h356 == io_rdAddr_0 ? lvtReg_854 : _GEN_4949; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4951 = 10'h357 == io_rdAddr_0 ? lvtReg_855 : _GEN_4950; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4952 = 10'h358 == io_rdAddr_0 ? lvtReg_856 : _GEN_4951; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4953 = 10'h359 == io_rdAddr_0 ? lvtReg_857 : _GEN_4952; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4954 = 10'h35a == io_rdAddr_0 ? lvtReg_858 : _GEN_4953; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4955 = 10'h35b == io_rdAddr_0 ? lvtReg_859 : _GEN_4954; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4956 = 10'h35c == io_rdAddr_0 ? lvtReg_860 : _GEN_4955; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4957 = 10'h35d == io_rdAddr_0 ? lvtReg_861 : _GEN_4956; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4958 = 10'h35e == io_rdAddr_0 ? lvtReg_862 : _GEN_4957; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4959 = 10'h35f == io_rdAddr_0 ? lvtReg_863 : _GEN_4958; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4960 = 10'h360 == io_rdAddr_0 ? lvtReg_864 : _GEN_4959; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4961 = 10'h361 == io_rdAddr_0 ? lvtReg_865 : _GEN_4960; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4962 = 10'h362 == io_rdAddr_0 ? lvtReg_866 : _GEN_4961; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4963 = 10'h363 == io_rdAddr_0 ? lvtReg_867 : _GEN_4962; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4964 = 10'h364 == io_rdAddr_0 ? lvtReg_868 : _GEN_4963; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4965 = 10'h365 == io_rdAddr_0 ? lvtReg_869 : _GEN_4964; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4966 = 10'h366 == io_rdAddr_0 ? lvtReg_870 : _GEN_4965; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4967 = 10'h367 == io_rdAddr_0 ? lvtReg_871 : _GEN_4966; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4968 = 10'h368 == io_rdAddr_0 ? lvtReg_872 : _GEN_4967; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4969 = 10'h369 == io_rdAddr_0 ? lvtReg_873 : _GEN_4968; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4970 = 10'h36a == io_rdAddr_0 ? lvtReg_874 : _GEN_4969; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4971 = 10'h36b == io_rdAddr_0 ? lvtReg_875 : _GEN_4970; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4972 = 10'h36c == io_rdAddr_0 ? lvtReg_876 : _GEN_4971; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4973 = 10'h36d == io_rdAddr_0 ? lvtReg_877 : _GEN_4972; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4974 = 10'h36e == io_rdAddr_0 ? lvtReg_878 : _GEN_4973; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4975 = 10'h36f == io_rdAddr_0 ? lvtReg_879 : _GEN_4974; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4976 = 10'h370 == io_rdAddr_0 ? lvtReg_880 : _GEN_4975; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4977 = 10'h371 == io_rdAddr_0 ? lvtReg_881 : _GEN_4976; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4978 = 10'h372 == io_rdAddr_0 ? lvtReg_882 : _GEN_4977; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4979 = 10'h373 == io_rdAddr_0 ? lvtReg_883 : _GEN_4978; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4980 = 10'h374 == io_rdAddr_0 ? lvtReg_884 : _GEN_4979; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4981 = 10'h375 == io_rdAddr_0 ? lvtReg_885 : _GEN_4980; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4982 = 10'h376 == io_rdAddr_0 ? lvtReg_886 : _GEN_4981; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4983 = 10'h377 == io_rdAddr_0 ? lvtReg_887 : _GEN_4982; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4984 = 10'h378 == io_rdAddr_0 ? lvtReg_888 : _GEN_4983; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4985 = 10'h379 == io_rdAddr_0 ? lvtReg_889 : _GEN_4984; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4986 = 10'h37a == io_rdAddr_0 ? lvtReg_890 : _GEN_4985; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4987 = 10'h37b == io_rdAddr_0 ? lvtReg_891 : _GEN_4986; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4988 = 10'h37c == io_rdAddr_0 ? lvtReg_892 : _GEN_4987; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4989 = 10'h37d == io_rdAddr_0 ? lvtReg_893 : _GEN_4988; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4990 = 10'h37e == io_rdAddr_0 ? lvtReg_894 : _GEN_4989; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4991 = 10'h37f == io_rdAddr_0 ? lvtReg_895 : _GEN_4990; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4992 = 10'h380 == io_rdAddr_0 ? lvtReg_896 : _GEN_4991; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4993 = 10'h381 == io_rdAddr_0 ? lvtReg_897 : _GEN_4992; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4994 = 10'h382 == io_rdAddr_0 ? lvtReg_898 : _GEN_4993; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4995 = 10'h383 == io_rdAddr_0 ? lvtReg_899 : _GEN_4994; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4996 = 10'h384 == io_rdAddr_0 ? lvtReg_900 : _GEN_4995; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4997 = 10'h385 == io_rdAddr_0 ? lvtReg_901 : _GEN_4996; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4998 = 10'h386 == io_rdAddr_0 ? lvtReg_902 : _GEN_4997; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_4999 = 10'h387 == io_rdAddr_0 ? lvtReg_903 : _GEN_4998; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5000 = 10'h388 == io_rdAddr_0 ? lvtReg_904 : _GEN_4999; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5001 = 10'h389 == io_rdAddr_0 ? lvtReg_905 : _GEN_5000; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5002 = 10'h38a == io_rdAddr_0 ? lvtReg_906 : _GEN_5001; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5003 = 10'h38b == io_rdAddr_0 ? lvtReg_907 : _GEN_5002; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5004 = 10'h38c == io_rdAddr_0 ? lvtReg_908 : _GEN_5003; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5005 = 10'h38d == io_rdAddr_0 ? lvtReg_909 : _GEN_5004; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5006 = 10'h38e == io_rdAddr_0 ? lvtReg_910 : _GEN_5005; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5007 = 10'h38f == io_rdAddr_0 ? lvtReg_911 : _GEN_5006; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5008 = 10'h390 == io_rdAddr_0 ? lvtReg_912 : _GEN_5007; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5009 = 10'h391 == io_rdAddr_0 ? lvtReg_913 : _GEN_5008; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5010 = 10'h392 == io_rdAddr_0 ? lvtReg_914 : _GEN_5009; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5011 = 10'h393 == io_rdAddr_0 ? lvtReg_915 : _GEN_5010; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5012 = 10'h394 == io_rdAddr_0 ? lvtReg_916 : _GEN_5011; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5013 = 10'h395 == io_rdAddr_0 ? lvtReg_917 : _GEN_5012; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5014 = 10'h396 == io_rdAddr_0 ? lvtReg_918 : _GEN_5013; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5015 = 10'h397 == io_rdAddr_0 ? lvtReg_919 : _GEN_5014; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5016 = 10'h398 == io_rdAddr_0 ? lvtReg_920 : _GEN_5015; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5017 = 10'h399 == io_rdAddr_0 ? lvtReg_921 : _GEN_5016; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5018 = 10'h39a == io_rdAddr_0 ? lvtReg_922 : _GEN_5017; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5019 = 10'h39b == io_rdAddr_0 ? lvtReg_923 : _GEN_5018; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5020 = 10'h39c == io_rdAddr_0 ? lvtReg_924 : _GEN_5019; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5021 = 10'h39d == io_rdAddr_0 ? lvtReg_925 : _GEN_5020; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5022 = 10'h39e == io_rdAddr_0 ? lvtReg_926 : _GEN_5021; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5023 = 10'h39f == io_rdAddr_0 ? lvtReg_927 : _GEN_5022; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5024 = 10'h3a0 == io_rdAddr_0 ? lvtReg_928 : _GEN_5023; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5025 = 10'h3a1 == io_rdAddr_0 ? lvtReg_929 : _GEN_5024; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5026 = 10'h3a2 == io_rdAddr_0 ? lvtReg_930 : _GEN_5025; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5027 = 10'h3a3 == io_rdAddr_0 ? lvtReg_931 : _GEN_5026; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5028 = 10'h3a4 == io_rdAddr_0 ? lvtReg_932 : _GEN_5027; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5029 = 10'h3a5 == io_rdAddr_0 ? lvtReg_933 : _GEN_5028; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5030 = 10'h3a6 == io_rdAddr_0 ? lvtReg_934 : _GEN_5029; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5031 = 10'h3a7 == io_rdAddr_0 ? lvtReg_935 : _GEN_5030; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5032 = 10'h3a8 == io_rdAddr_0 ? lvtReg_936 : _GEN_5031; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5033 = 10'h3a9 == io_rdAddr_0 ? lvtReg_937 : _GEN_5032; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5034 = 10'h3aa == io_rdAddr_0 ? lvtReg_938 : _GEN_5033; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5035 = 10'h3ab == io_rdAddr_0 ? lvtReg_939 : _GEN_5034; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5036 = 10'h3ac == io_rdAddr_0 ? lvtReg_940 : _GEN_5035; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5037 = 10'h3ad == io_rdAddr_0 ? lvtReg_941 : _GEN_5036; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5038 = 10'h3ae == io_rdAddr_0 ? lvtReg_942 : _GEN_5037; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5039 = 10'h3af == io_rdAddr_0 ? lvtReg_943 : _GEN_5038; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5040 = 10'h3b0 == io_rdAddr_0 ? lvtReg_944 : _GEN_5039; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5041 = 10'h3b1 == io_rdAddr_0 ? lvtReg_945 : _GEN_5040; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5042 = 10'h3b2 == io_rdAddr_0 ? lvtReg_946 : _GEN_5041; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5043 = 10'h3b3 == io_rdAddr_0 ? lvtReg_947 : _GEN_5042; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5044 = 10'h3b4 == io_rdAddr_0 ? lvtReg_948 : _GEN_5043; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5045 = 10'h3b5 == io_rdAddr_0 ? lvtReg_949 : _GEN_5044; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5046 = 10'h3b6 == io_rdAddr_0 ? lvtReg_950 : _GEN_5045; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5047 = 10'h3b7 == io_rdAddr_0 ? lvtReg_951 : _GEN_5046; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5048 = 10'h3b8 == io_rdAddr_0 ? lvtReg_952 : _GEN_5047; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5049 = 10'h3b9 == io_rdAddr_0 ? lvtReg_953 : _GEN_5048; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5050 = 10'h3ba == io_rdAddr_0 ? lvtReg_954 : _GEN_5049; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5051 = 10'h3bb == io_rdAddr_0 ? lvtReg_955 : _GEN_5050; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5052 = 10'h3bc == io_rdAddr_0 ? lvtReg_956 : _GEN_5051; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5053 = 10'h3bd == io_rdAddr_0 ? lvtReg_957 : _GEN_5052; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5054 = 10'h3be == io_rdAddr_0 ? lvtReg_958 : _GEN_5053; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5055 = 10'h3bf == io_rdAddr_0 ? lvtReg_959 : _GEN_5054; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5056 = 10'h3c0 == io_rdAddr_0 ? lvtReg_960 : _GEN_5055; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5057 = 10'h3c1 == io_rdAddr_0 ? lvtReg_961 : _GEN_5056; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5058 = 10'h3c2 == io_rdAddr_0 ? lvtReg_962 : _GEN_5057; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5059 = 10'h3c3 == io_rdAddr_0 ? lvtReg_963 : _GEN_5058; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5060 = 10'h3c4 == io_rdAddr_0 ? lvtReg_964 : _GEN_5059; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5061 = 10'h3c5 == io_rdAddr_0 ? lvtReg_965 : _GEN_5060; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5062 = 10'h3c6 == io_rdAddr_0 ? lvtReg_966 : _GEN_5061; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5063 = 10'h3c7 == io_rdAddr_0 ? lvtReg_967 : _GEN_5062; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5064 = 10'h3c8 == io_rdAddr_0 ? lvtReg_968 : _GEN_5063; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5065 = 10'h3c9 == io_rdAddr_0 ? lvtReg_969 : _GEN_5064; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5066 = 10'h3ca == io_rdAddr_0 ? lvtReg_970 : _GEN_5065; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5067 = 10'h3cb == io_rdAddr_0 ? lvtReg_971 : _GEN_5066; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5068 = 10'h3cc == io_rdAddr_0 ? lvtReg_972 : _GEN_5067; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5069 = 10'h3cd == io_rdAddr_0 ? lvtReg_973 : _GEN_5068; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5070 = 10'h3ce == io_rdAddr_0 ? lvtReg_974 : _GEN_5069; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5071 = 10'h3cf == io_rdAddr_0 ? lvtReg_975 : _GEN_5070; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5072 = 10'h3d0 == io_rdAddr_0 ? lvtReg_976 : _GEN_5071; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5073 = 10'h3d1 == io_rdAddr_0 ? lvtReg_977 : _GEN_5072; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5074 = 10'h3d2 == io_rdAddr_0 ? lvtReg_978 : _GEN_5073; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5075 = 10'h3d3 == io_rdAddr_0 ? lvtReg_979 : _GEN_5074; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5076 = 10'h3d4 == io_rdAddr_0 ? lvtReg_980 : _GEN_5075; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5077 = 10'h3d5 == io_rdAddr_0 ? lvtReg_981 : _GEN_5076; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5078 = 10'h3d6 == io_rdAddr_0 ? lvtReg_982 : _GEN_5077; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5079 = 10'h3d7 == io_rdAddr_0 ? lvtReg_983 : _GEN_5078; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5080 = 10'h3d8 == io_rdAddr_0 ? lvtReg_984 : _GEN_5079; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5081 = 10'h3d9 == io_rdAddr_0 ? lvtReg_985 : _GEN_5080; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5082 = 10'h3da == io_rdAddr_0 ? lvtReg_986 : _GEN_5081; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5083 = 10'h3db == io_rdAddr_0 ? lvtReg_987 : _GEN_5082; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5084 = 10'h3dc == io_rdAddr_0 ? lvtReg_988 : _GEN_5083; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5085 = 10'h3dd == io_rdAddr_0 ? lvtReg_989 : _GEN_5084; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5086 = 10'h3de == io_rdAddr_0 ? lvtReg_990 : _GEN_5085; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5087 = 10'h3df == io_rdAddr_0 ? lvtReg_991 : _GEN_5086; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5088 = 10'h3e0 == io_rdAddr_0 ? lvtReg_992 : _GEN_5087; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5089 = 10'h3e1 == io_rdAddr_0 ? lvtReg_993 : _GEN_5088; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5090 = 10'h3e2 == io_rdAddr_0 ? lvtReg_994 : _GEN_5089; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5091 = 10'h3e3 == io_rdAddr_0 ? lvtReg_995 : _GEN_5090; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5092 = 10'h3e4 == io_rdAddr_0 ? lvtReg_996 : _GEN_5091; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5093 = 10'h3e5 == io_rdAddr_0 ? lvtReg_997 : _GEN_5092; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5094 = 10'h3e6 == io_rdAddr_0 ? lvtReg_998 : _GEN_5093; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5095 = 10'h3e7 == io_rdAddr_0 ? lvtReg_999 : _GEN_5094; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5096 = 10'h3e8 == io_rdAddr_0 ? lvtReg_1000 : _GEN_5095; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5097 = 10'h3e9 == io_rdAddr_0 ? lvtReg_1001 : _GEN_5096; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5098 = 10'h3ea == io_rdAddr_0 ? lvtReg_1002 : _GEN_5097; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5099 = 10'h3eb == io_rdAddr_0 ? lvtReg_1003 : _GEN_5098; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5100 = 10'h3ec == io_rdAddr_0 ? lvtReg_1004 : _GEN_5099; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5101 = 10'h3ed == io_rdAddr_0 ? lvtReg_1005 : _GEN_5100; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5102 = 10'h3ee == io_rdAddr_0 ? lvtReg_1006 : _GEN_5101; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5103 = 10'h3ef == io_rdAddr_0 ? lvtReg_1007 : _GEN_5102; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5104 = 10'h3f0 == io_rdAddr_0 ? lvtReg_1008 : _GEN_5103; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5105 = 10'h3f1 == io_rdAddr_0 ? lvtReg_1009 : _GEN_5104; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5106 = 10'h3f2 == io_rdAddr_0 ? lvtReg_1010 : _GEN_5105; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5107 = 10'h3f3 == io_rdAddr_0 ? lvtReg_1011 : _GEN_5106; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5108 = 10'h3f4 == io_rdAddr_0 ? lvtReg_1012 : _GEN_5107; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5109 = 10'h3f5 == io_rdAddr_0 ? lvtReg_1013 : _GEN_5108; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5110 = 10'h3f6 == io_rdAddr_0 ? lvtReg_1014 : _GEN_5109; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5111 = 10'h3f7 == io_rdAddr_0 ? lvtReg_1015 : _GEN_5110; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5112 = 10'h3f8 == io_rdAddr_0 ? lvtReg_1016 : _GEN_5111; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5113 = 10'h3f9 == io_rdAddr_0 ? lvtReg_1017 : _GEN_5112; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5114 = 10'h3fa == io_rdAddr_0 ? lvtReg_1018 : _GEN_5113; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5115 = 10'h3fb == io_rdAddr_0 ? lvtReg_1019 : _GEN_5114; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5116 = 10'h3fc == io_rdAddr_0 ? lvtReg_1020 : _GEN_5115; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5117 = 10'h3fd == io_rdAddr_0 ? lvtReg_1021 : _GEN_5116; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5118 = 10'h3fe == io_rdAddr_0 ? lvtReg_1022 : _GEN_5117; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5121 = 10'h1 == io_rdAddr_1 ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5122 = 10'h2 == io_rdAddr_1 ? lvtReg_2 : _GEN_5121; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5123 = 10'h3 == io_rdAddr_1 ? lvtReg_3 : _GEN_5122; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5124 = 10'h4 == io_rdAddr_1 ? lvtReg_4 : _GEN_5123; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5125 = 10'h5 == io_rdAddr_1 ? lvtReg_5 : _GEN_5124; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5126 = 10'h6 == io_rdAddr_1 ? lvtReg_6 : _GEN_5125; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5127 = 10'h7 == io_rdAddr_1 ? lvtReg_7 : _GEN_5126; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5128 = 10'h8 == io_rdAddr_1 ? lvtReg_8 : _GEN_5127; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5129 = 10'h9 == io_rdAddr_1 ? lvtReg_9 : _GEN_5128; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5130 = 10'ha == io_rdAddr_1 ? lvtReg_10 : _GEN_5129; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5131 = 10'hb == io_rdAddr_1 ? lvtReg_11 : _GEN_5130; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5132 = 10'hc == io_rdAddr_1 ? lvtReg_12 : _GEN_5131; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5133 = 10'hd == io_rdAddr_1 ? lvtReg_13 : _GEN_5132; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5134 = 10'he == io_rdAddr_1 ? lvtReg_14 : _GEN_5133; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5135 = 10'hf == io_rdAddr_1 ? lvtReg_15 : _GEN_5134; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5136 = 10'h10 == io_rdAddr_1 ? lvtReg_16 : _GEN_5135; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5137 = 10'h11 == io_rdAddr_1 ? lvtReg_17 : _GEN_5136; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5138 = 10'h12 == io_rdAddr_1 ? lvtReg_18 : _GEN_5137; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5139 = 10'h13 == io_rdAddr_1 ? lvtReg_19 : _GEN_5138; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5140 = 10'h14 == io_rdAddr_1 ? lvtReg_20 : _GEN_5139; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5141 = 10'h15 == io_rdAddr_1 ? lvtReg_21 : _GEN_5140; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5142 = 10'h16 == io_rdAddr_1 ? lvtReg_22 : _GEN_5141; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5143 = 10'h17 == io_rdAddr_1 ? lvtReg_23 : _GEN_5142; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5144 = 10'h18 == io_rdAddr_1 ? lvtReg_24 : _GEN_5143; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5145 = 10'h19 == io_rdAddr_1 ? lvtReg_25 : _GEN_5144; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5146 = 10'h1a == io_rdAddr_1 ? lvtReg_26 : _GEN_5145; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5147 = 10'h1b == io_rdAddr_1 ? lvtReg_27 : _GEN_5146; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5148 = 10'h1c == io_rdAddr_1 ? lvtReg_28 : _GEN_5147; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5149 = 10'h1d == io_rdAddr_1 ? lvtReg_29 : _GEN_5148; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5150 = 10'h1e == io_rdAddr_1 ? lvtReg_30 : _GEN_5149; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5151 = 10'h1f == io_rdAddr_1 ? lvtReg_31 : _GEN_5150; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5152 = 10'h20 == io_rdAddr_1 ? lvtReg_32 : _GEN_5151; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5153 = 10'h21 == io_rdAddr_1 ? lvtReg_33 : _GEN_5152; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5154 = 10'h22 == io_rdAddr_1 ? lvtReg_34 : _GEN_5153; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5155 = 10'h23 == io_rdAddr_1 ? lvtReg_35 : _GEN_5154; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5156 = 10'h24 == io_rdAddr_1 ? lvtReg_36 : _GEN_5155; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5157 = 10'h25 == io_rdAddr_1 ? lvtReg_37 : _GEN_5156; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5158 = 10'h26 == io_rdAddr_1 ? lvtReg_38 : _GEN_5157; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5159 = 10'h27 == io_rdAddr_1 ? lvtReg_39 : _GEN_5158; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5160 = 10'h28 == io_rdAddr_1 ? lvtReg_40 : _GEN_5159; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5161 = 10'h29 == io_rdAddr_1 ? lvtReg_41 : _GEN_5160; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5162 = 10'h2a == io_rdAddr_1 ? lvtReg_42 : _GEN_5161; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5163 = 10'h2b == io_rdAddr_1 ? lvtReg_43 : _GEN_5162; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5164 = 10'h2c == io_rdAddr_1 ? lvtReg_44 : _GEN_5163; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5165 = 10'h2d == io_rdAddr_1 ? lvtReg_45 : _GEN_5164; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5166 = 10'h2e == io_rdAddr_1 ? lvtReg_46 : _GEN_5165; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5167 = 10'h2f == io_rdAddr_1 ? lvtReg_47 : _GEN_5166; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5168 = 10'h30 == io_rdAddr_1 ? lvtReg_48 : _GEN_5167; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5169 = 10'h31 == io_rdAddr_1 ? lvtReg_49 : _GEN_5168; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5170 = 10'h32 == io_rdAddr_1 ? lvtReg_50 : _GEN_5169; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5171 = 10'h33 == io_rdAddr_1 ? lvtReg_51 : _GEN_5170; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5172 = 10'h34 == io_rdAddr_1 ? lvtReg_52 : _GEN_5171; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5173 = 10'h35 == io_rdAddr_1 ? lvtReg_53 : _GEN_5172; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5174 = 10'h36 == io_rdAddr_1 ? lvtReg_54 : _GEN_5173; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5175 = 10'h37 == io_rdAddr_1 ? lvtReg_55 : _GEN_5174; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5176 = 10'h38 == io_rdAddr_1 ? lvtReg_56 : _GEN_5175; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5177 = 10'h39 == io_rdAddr_1 ? lvtReg_57 : _GEN_5176; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5178 = 10'h3a == io_rdAddr_1 ? lvtReg_58 : _GEN_5177; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5179 = 10'h3b == io_rdAddr_1 ? lvtReg_59 : _GEN_5178; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5180 = 10'h3c == io_rdAddr_1 ? lvtReg_60 : _GEN_5179; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5181 = 10'h3d == io_rdAddr_1 ? lvtReg_61 : _GEN_5180; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5182 = 10'h3e == io_rdAddr_1 ? lvtReg_62 : _GEN_5181; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5183 = 10'h3f == io_rdAddr_1 ? lvtReg_63 : _GEN_5182; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5184 = 10'h40 == io_rdAddr_1 ? lvtReg_64 : _GEN_5183; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5185 = 10'h41 == io_rdAddr_1 ? lvtReg_65 : _GEN_5184; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5186 = 10'h42 == io_rdAddr_1 ? lvtReg_66 : _GEN_5185; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5187 = 10'h43 == io_rdAddr_1 ? lvtReg_67 : _GEN_5186; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5188 = 10'h44 == io_rdAddr_1 ? lvtReg_68 : _GEN_5187; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5189 = 10'h45 == io_rdAddr_1 ? lvtReg_69 : _GEN_5188; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5190 = 10'h46 == io_rdAddr_1 ? lvtReg_70 : _GEN_5189; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5191 = 10'h47 == io_rdAddr_1 ? lvtReg_71 : _GEN_5190; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5192 = 10'h48 == io_rdAddr_1 ? lvtReg_72 : _GEN_5191; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5193 = 10'h49 == io_rdAddr_1 ? lvtReg_73 : _GEN_5192; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5194 = 10'h4a == io_rdAddr_1 ? lvtReg_74 : _GEN_5193; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5195 = 10'h4b == io_rdAddr_1 ? lvtReg_75 : _GEN_5194; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5196 = 10'h4c == io_rdAddr_1 ? lvtReg_76 : _GEN_5195; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5197 = 10'h4d == io_rdAddr_1 ? lvtReg_77 : _GEN_5196; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5198 = 10'h4e == io_rdAddr_1 ? lvtReg_78 : _GEN_5197; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5199 = 10'h4f == io_rdAddr_1 ? lvtReg_79 : _GEN_5198; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5200 = 10'h50 == io_rdAddr_1 ? lvtReg_80 : _GEN_5199; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5201 = 10'h51 == io_rdAddr_1 ? lvtReg_81 : _GEN_5200; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5202 = 10'h52 == io_rdAddr_1 ? lvtReg_82 : _GEN_5201; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5203 = 10'h53 == io_rdAddr_1 ? lvtReg_83 : _GEN_5202; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5204 = 10'h54 == io_rdAddr_1 ? lvtReg_84 : _GEN_5203; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5205 = 10'h55 == io_rdAddr_1 ? lvtReg_85 : _GEN_5204; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5206 = 10'h56 == io_rdAddr_1 ? lvtReg_86 : _GEN_5205; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5207 = 10'h57 == io_rdAddr_1 ? lvtReg_87 : _GEN_5206; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5208 = 10'h58 == io_rdAddr_1 ? lvtReg_88 : _GEN_5207; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5209 = 10'h59 == io_rdAddr_1 ? lvtReg_89 : _GEN_5208; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5210 = 10'h5a == io_rdAddr_1 ? lvtReg_90 : _GEN_5209; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5211 = 10'h5b == io_rdAddr_1 ? lvtReg_91 : _GEN_5210; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5212 = 10'h5c == io_rdAddr_1 ? lvtReg_92 : _GEN_5211; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5213 = 10'h5d == io_rdAddr_1 ? lvtReg_93 : _GEN_5212; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5214 = 10'h5e == io_rdAddr_1 ? lvtReg_94 : _GEN_5213; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5215 = 10'h5f == io_rdAddr_1 ? lvtReg_95 : _GEN_5214; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5216 = 10'h60 == io_rdAddr_1 ? lvtReg_96 : _GEN_5215; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5217 = 10'h61 == io_rdAddr_1 ? lvtReg_97 : _GEN_5216; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5218 = 10'h62 == io_rdAddr_1 ? lvtReg_98 : _GEN_5217; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5219 = 10'h63 == io_rdAddr_1 ? lvtReg_99 : _GEN_5218; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5220 = 10'h64 == io_rdAddr_1 ? lvtReg_100 : _GEN_5219; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5221 = 10'h65 == io_rdAddr_1 ? lvtReg_101 : _GEN_5220; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5222 = 10'h66 == io_rdAddr_1 ? lvtReg_102 : _GEN_5221; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5223 = 10'h67 == io_rdAddr_1 ? lvtReg_103 : _GEN_5222; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5224 = 10'h68 == io_rdAddr_1 ? lvtReg_104 : _GEN_5223; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5225 = 10'h69 == io_rdAddr_1 ? lvtReg_105 : _GEN_5224; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5226 = 10'h6a == io_rdAddr_1 ? lvtReg_106 : _GEN_5225; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5227 = 10'h6b == io_rdAddr_1 ? lvtReg_107 : _GEN_5226; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5228 = 10'h6c == io_rdAddr_1 ? lvtReg_108 : _GEN_5227; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5229 = 10'h6d == io_rdAddr_1 ? lvtReg_109 : _GEN_5228; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5230 = 10'h6e == io_rdAddr_1 ? lvtReg_110 : _GEN_5229; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5231 = 10'h6f == io_rdAddr_1 ? lvtReg_111 : _GEN_5230; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5232 = 10'h70 == io_rdAddr_1 ? lvtReg_112 : _GEN_5231; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5233 = 10'h71 == io_rdAddr_1 ? lvtReg_113 : _GEN_5232; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5234 = 10'h72 == io_rdAddr_1 ? lvtReg_114 : _GEN_5233; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5235 = 10'h73 == io_rdAddr_1 ? lvtReg_115 : _GEN_5234; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5236 = 10'h74 == io_rdAddr_1 ? lvtReg_116 : _GEN_5235; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5237 = 10'h75 == io_rdAddr_1 ? lvtReg_117 : _GEN_5236; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5238 = 10'h76 == io_rdAddr_1 ? lvtReg_118 : _GEN_5237; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5239 = 10'h77 == io_rdAddr_1 ? lvtReg_119 : _GEN_5238; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5240 = 10'h78 == io_rdAddr_1 ? lvtReg_120 : _GEN_5239; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5241 = 10'h79 == io_rdAddr_1 ? lvtReg_121 : _GEN_5240; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5242 = 10'h7a == io_rdAddr_1 ? lvtReg_122 : _GEN_5241; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5243 = 10'h7b == io_rdAddr_1 ? lvtReg_123 : _GEN_5242; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5244 = 10'h7c == io_rdAddr_1 ? lvtReg_124 : _GEN_5243; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5245 = 10'h7d == io_rdAddr_1 ? lvtReg_125 : _GEN_5244; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5246 = 10'h7e == io_rdAddr_1 ? lvtReg_126 : _GEN_5245; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5247 = 10'h7f == io_rdAddr_1 ? lvtReg_127 : _GEN_5246; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5248 = 10'h80 == io_rdAddr_1 ? lvtReg_128 : _GEN_5247; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5249 = 10'h81 == io_rdAddr_1 ? lvtReg_129 : _GEN_5248; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5250 = 10'h82 == io_rdAddr_1 ? lvtReg_130 : _GEN_5249; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5251 = 10'h83 == io_rdAddr_1 ? lvtReg_131 : _GEN_5250; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5252 = 10'h84 == io_rdAddr_1 ? lvtReg_132 : _GEN_5251; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5253 = 10'h85 == io_rdAddr_1 ? lvtReg_133 : _GEN_5252; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5254 = 10'h86 == io_rdAddr_1 ? lvtReg_134 : _GEN_5253; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5255 = 10'h87 == io_rdAddr_1 ? lvtReg_135 : _GEN_5254; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5256 = 10'h88 == io_rdAddr_1 ? lvtReg_136 : _GEN_5255; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5257 = 10'h89 == io_rdAddr_1 ? lvtReg_137 : _GEN_5256; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5258 = 10'h8a == io_rdAddr_1 ? lvtReg_138 : _GEN_5257; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5259 = 10'h8b == io_rdAddr_1 ? lvtReg_139 : _GEN_5258; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5260 = 10'h8c == io_rdAddr_1 ? lvtReg_140 : _GEN_5259; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5261 = 10'h8d == io_rdAddr_1 ? lvtReg_141 : _GEN_5260; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5262 = 10'h8e == io_rdAddr_1 ? lvtReg_142 : _GEN_5261; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5263 = 10'h8f == io_rdAddr_1 ? lvtReg_143 : _GEN_5262; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5264 = 10'h90 == io_rdAddr_1 ? lvtReg_144 : _GEN_5263; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5265 = 10'h91 == io_rdAddr_1 ? lvtReg_145 : _GEN_5264; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5266 = 10'h92 == io_rdAddr_1 ? lvtReg_146 : _GEN_5265; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5267 = 10'h93 == io_rdAddr_1 ? lvtReg_147 : _GEN_5266; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5268 = 10'h94 == io_rdAddr_1 ? lvtReg_148 : _GEN_5267; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5269 = 10'h95 == io_rdAddr_1 ? lvtReg_149 : _GEN_5268; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5270 = 10'h96 == io_rdAddr_1 ? lvtReg_150 : _GEN_5269; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5271 = 10'h97 == io_rdAddr_1 ? lvtReg_151 : _GEN_5270; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5272 = 10'h98 == io_rdAddr_1 ? lvtReg_152 : _GEN_5271; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5273 = 10'h99 == io_rdAddr_1 ? lvtReg_153 : _GEN_5272; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5274 = 10'h9a == io_rdAddr_1 ? lvtReg_154 : _GEN_5273; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5275 = 10'h9b == io_rdAddr_1 ? lvtReg_155 : _GEN_5274; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5276 = 10'h9c == io_rdAddr_1 ? lvtReg_156 : _GEN_5275; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5277 = 10'h9d == io_rdAddr_1 ? lvtReg_157 : _GEN_5276; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5278 = 10'h9e == io_rdAddr_1 ? lvtReg_158 : _GEN_5277; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5279 = 10'h9f == io_rdAddr_1 ? lvtReg_159 : _GEN_5278; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5280 = 10'ha0 == io_rdAddr_1 ? lvtReg_160 : _GEN_5279; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5281 = 10'ha1 == io_rdAddr_1 ? lvtReg_161 : _GEN_5280; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5282 = 10'ha2 == io_rdAddr_1 ? lvtReg_162 : _GEN_5281; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5283 = 10'ha3 == io_rdAddr_1 ? lvtReg_163 : _GEN_5282; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5284 = 10'ha4 == io_rdAddr_1 ? lvtReg_164 : _GEN_5283; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5285 = 10'ha5 == io_rdAddr_1 ? lvtReg_165 : _GEN_5284; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5286 = 10'ha6 == io_rdAddr_1 ? lvtReg_166 : _GEN_5285; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5287 = 10'ha7 == io_rdAddr_1 ? lvtReg_167 : _GEN_5286; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5288 = 10'ha8 == io_rdAddr_1 ? lvtReg_168 : _GEN_5287; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5289 = 10'ha9 == io_rdAddr_1 ? lvtReg_169 : _GEN_5288; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5290 = 10'haa == io_rdAddr_1 ? lvtReg_170 : _GEN_5289; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5291 = 10'hab == io_rdAddr_1 ? lvtReg_171 : _GEN_5290; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5292 = 10'hac == io_rdAddr_1 ? lvtReg_172 : _GEN_5291; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5293 = 10'had == io_rdAddr_1 ? lvtReg_173 : _GEN_5292; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5294 = 10'hae == io_rdAddr_1 ? lvtReg_174 : _GEN_5293; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5295 = 10'haf == io_rdAddr_1 ? lvtReg_175 : _GEN_5294; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5296 = 10'hb0 == io_rdAddr_1 ? lvtReg_176 : _GEN_5295; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5297 = 10'hb1 == io_rdAddr_1 ? lvtReg_177 : _GEN_5296; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5298 = 10'hb2 == io_rdAddr_1 ? lvtReg_178 : _GEN_5297; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5299 = 10'hb3 == io_rdAddr_1 ? lvtReg_179 : _GEN_5298; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5300 = 10'hb4 == io_rdAddr_1 ? lvtReg_180 : _GEN_5299; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5301 = 10'hb5 == io_rdAddr_1 ? lvtReg_181 : _GEN_5300; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5302 = 10'hb6 == io_rdAddr_1 ? lvtReg_182 : _GEN_5301; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5303 = 10'hb7 == io_rdAddr_1 ? lvtReg_183 : _GEN_5302; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5304 = 10'hb8 == io_rdAddr_1 ? lvtReg_184 : _GEN_5303; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5305 = 10'hb9 == io_rdAddr_1 ? lvtReg_185 : _GEN_5304; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5306 = 10'hba == io_rdAddr_1 ? lvtReg_186 : _GEN_5305; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5307 = 10'hbb == io_rdAddr_1 ? lvtReg_187 : _GEN_5306; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5308 = 10'hbc == io_rdAddr_1 ? lvtReg_188 : _GEN_5307; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5309 = 10'hbd == io_rdAddr_1 ? lvtReg_189 : _GEN_5308; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5310 = 10'hbe == io_rdAddr_1 ? lvtReg_190 : _GEN_5309; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5311 = 10'hbf == io_rdAddr_1 ? lvtReg_191 : _GEN_5310; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5312 = 10'hc0 == io_rdAddr_1 ? lvtReg_192 : _GEN_5311; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5313 = 10'hc1 == io_rdAddr_1 ? lvtReg_193 : _GEN_5312; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5314 = 10'hc2 == io_rdAddr_1 ? lvtReg_194 : _GEN_5313; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5315 = 10'hc3 == io_rdAddr_1 ? lvtReg_195 : _GEN_5314; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5316 = 10'hc4 == io_rdAddr_1 ? lvtReg_196 : _GEN_5315; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5317 = 10'hc5 == io_rdAddr_1 ? lvtReg_197 : _GEN_5316; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5318 = 10'hc6 == io_rdAddr_1 ? lvtReg_198 : _GEN_5317; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5319 = 10'hc7 == io_rdAddr_1 ? lvtReg_199 : _GEN_5318; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5320 = 10'hc8 == io_rdAddr_1 ? lvtReg_200 : _GEN_5319; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5321 = 10'hc9 == io_rdAddr_1 ? lvtReg_201 : _GEN_5320; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5322 = 10'hca == io_rdAddr_1 ? lvtReg_202 : _GEN_5321; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5323 = 10'hcb == io_rdAddr_1 ? lvtReg_203 : _GEN_5322; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5324 = 10'hcc == io_rdAddr_1 ? lvtReg_204 : _GEN_5323; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5325 = 10'hcd == io_rdAddr_1 ? lvtReg_205 : _GEN_5324; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5326 = 10'hce == io_rdAddr_1 ? lvtReg_206 : _GEN_5325; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5327 = 10'hcf == io_rdAddr_1 ? lvtReg_207 : _GEN_5326; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5328 = 10'hd0 == io_rdAddr_1 ? lvtReg_208 : _GEN_5327; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5329 = 10'hd1 == io_rdAddr_1 ? lvtReg_209 : _GEN_5328; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5330 = 10'hd2 == io_rdAddr_1 ? lvtReg_210 : _GEN_5329; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5331 = 10'hd3 == io_rdAddr_1 ? lvtReg_211 : _GEN_5330; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5332 = 10'hd4 == io_rdAddr_1 ? lvtReg_212 : _GEN_5331; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5333 = 10'hd5 == io_rdAddr_1 ? lvtReg_213 : _GEN_5332; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5334 = 10'hd6 == io_rdAddr_1 ? lvtReg_214 : _GEN_5333; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5335 = 10'hd7 == io_rdAddr_1 ? lvtReg_215 : _GEN_5334; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5336 = 10'hd8 == io_rdAddr_1 ? lvtReg_216 : _GEN_5335; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5337 = 10'hd9 == io_rdAddr_1 ? lvtReg_217 : _GEN_5336; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5338 = 10'hda == io_rdAddr_1 ? lvtReg_218 : _GEN_5337; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5339 = 10'hdb == io_rdAddr_1 ? lvtReg_219 : _GEN_5338; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5340 = 10'hdc == io_rdAddr_1 ? lvtReg_220 : _GEN_5339; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5341 = 10'hdd == io_rdAddr_1 ? lvtReg_221 : _GEN_5340; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5342 = 10'hde == io_rdAddr_1 ? lvtReg_222 : _GEN_5341; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5343 = 10'hdf == io_rdAddr_1 ? lvtReg_223 : _GEN_5342; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5344 = 10'he0 == io_rdAddr_1 ? lvtReg_224 : _GEN_5343; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5345 = 10'he1 == io_rdAddr_1 ? lvtReg_225 : _GEN_5344; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5346 = 10'he2 == io_rdAddr_1 ? lvtReg_226 : _GEN_5345; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5347 = 10'he3 == io_rdAddr_1 ? lvtReg_227 : _GEN_5346; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5348 = 10'he4 == io_rdAddr_1 ? lvtReg_228 : _GEN_5347; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5349 = 10'he5 == io_rdAddr_1 ? lvtReg_229 : _GEN_5348; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5350 = 10'he6 == io_rdAddr_1 ? lvtReg_230 : _GEN_5349; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5351 = 10'he7 == io_rdAddr_1 ? lvtReg_231 : _GEN_5350; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5352 = 10'he8 == io_rdAddr_1 ? lvtReg_232 : _GEN_5351; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5353 = 10'he9 == io_rdAddr_1 ? lvtReg_233 : _GEN_5352; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5354 = 10'hea == io_rdAddr_1 ? lvtReg_234 : _GEN_5353; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5355 = 10'heb == io_rdAddr_1 ? lvtReg_235 : _GEN_5354; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5356 = 10'hec == io_rdAddr_1 ? lvtReg_236 : _GEN_5355; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5357 = 10'hed == io_rdAddr_1 ? lvtReg_237 : _GEN_5356; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5358 = 10'hee == io_rdAddr_1 ? lvtReg_238 : _GEN_5357; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5359 = 10'hef == io_rdAddr_1 ? lvtReg_239 : _GEN_5358; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5360 = 10'hf0 == io_rdAddr_1 ? lvtReg_240 : _GEN_5359; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5361 = 10'hf1 == io_rdAddr_1 ? lvtReg_241 : _GEN_5360; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5362 = 10'hf2 == io_rdAddr_1 ? lvtReg_242 : _GEN_5361; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5363 = 10'hf3 == io_rdAddr_1 ? lvtReg_243 : _GEN_5362; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5364 = 10'hf4 == io_rdAddr_1 ? lvtReg_244 : _GEN_5363; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5365 = 10'hf5 == io_rdAddr_1 ? lvtReg_245 : _GEN_5364; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5366 = 10'hf6 == io_rdAddr_1 ? lvtReg_246 : _GEN_5365; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5367 = 10'hf7 == io_rdAddr_1 ? lvtReg_247 : _GEN_5366; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5368 = 10'hf8 == io_rdAddr_1 ? lvtReg_248 : _GEN_5367; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5369 = 10'hf9 == io_rdAddr_1 ? lvtReg_249 : _GEN_5368; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5370 = 10'hfa == io_rdAddr_1 ? lvtReg_250 : _GEN_5369; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5371 = 10'hfb == io_rdAddr_1 ? lvtReg_251 : _GEN_5370; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5372 = 10'hfc == io_rdAddr_1 ? lvtReg_252 : _GEN_5371; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5373 = 10'hfd == io_rdAddr_1 ? lvtReg_253 : _GEN_5372; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5374 = 10'hfe == io_rdAddr_1 ? lvtReg_254 : _GEN_5373; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5375 = 10'hff == io_rdAddr_1 ? lvtReg_255 : _GEN_5374; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5376 = 10'h100 == io_rdAddr_1 ? lvtReg_256 : _GEN_5375; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5377 = 10'h101 == io_rdAddr_1 ? lvtReg_257 : _GEN_5376; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5378 = 10'h102 == io_rdAddr_1 ? lvtReg_258 : _GEN_5377; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5379 = 10'h103 == io_rdAddr_1 ? lvtReg_259 : _GEN_5378; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5380 = 10'h104 == io_rdAddr_1 ? lvtReg_260 : _GEN_5379; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5381 = 10'h105 == io_rdAddr_1 ? lvtReg_261 : _GEN_5380; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5382 = 10'h106 == io_rdAddr_1 ? lvtReg_262 : _GEN_5381; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5383 = 10'h107 == io_rdAddr_1 ? lvtReg_263 : _GEN_5382; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5384 = 10'h108 == io_rdAddr_1 ? lvtReg_264 : _GEN_5383; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5385 = 10'h109 == io_rdAddr_1 ? lvtReg_265 : _GEN_5384; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5386 = 10'h10a == io_rdAddr_1 ? lvtReg_266 : _GEN_5385; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5387 = 10'h10b == io_rdAddr_1 ? lvtReg_267 : _GEN_5386; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5388 = 10'h10c == io_rdAddr_1 ? lvtReg_268 : _GEN_5387; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5389 = 10'h10d == io_rdAddr_1 ? lvtReg_269 : _GEN_5388; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5390 = 10'h10e == io_rdAddr_1 ? lvtReg_270 : _GEN_5389; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5391 = 10'h10f == io_rdAddr_1 ? lvtReg_271 : _GEN_5390; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5392 = 10'h110 == io_rdAddr_1 ? lvtReg_272 : _GEN_5391; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5393 = 10'h111 == io_rdAddr_1 ? lvtReg_273 : _GEN_5392; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5394 = 10'h112 == io_rdAddr_1 ? lvtReg_274 : _GEN_5393; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5395 = 10'h113 == io_rdAddr_1 ? lvtReg_275 : _GEN_5394; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5396 = 10'h114 == io_rdAddr_1 ? lvtReg_276 : _GEN_5395; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5397 = 10'h115 == io_rdAddr_1 ? lvtReg_277 : _GEN_5396; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5398 = 10'h116 == io_rdAddr_1 ? lvtReg_278 : _GEN_5397; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5399 = 10'h117 == io_rdAddr_1 ? lvtReg_279 : _GEN_5398; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5400 = 10'h118 == io_rdAddr_1 ? lvtReg_280 : _GEN_5399; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5401 = 10'h119 == io_rdAddr_1 ? lvtReg_281 : _GEN_5400; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5402 = 10'h11a == io_rdAddr_1 ? lvtReg_282 : _GEN_5401; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5403 = 10'h11b == io_rdAddr_1 ? lvtReg_283 : _GEN_5402; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5404 = 10'h11c == io_rdAddr_1 ? lvtReg_284 : _GEN_5403; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5405 = 10'h11d == io_rdAddr_1 ? lvtReg_285 : _GEN_5404; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5406 = 10'h11e == io_rdAddr_1 ? lvtReg_286 : _GEN_5405; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5407 = 10'h11f == io_rdAddr_1 ? lvtReg_287 : _GEN_5406; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5408 = 10'h120 == io_rdAddr_1 ? lvtReg_288 : _GEN_5407; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5409 = 10'h121 == io_rdAddr_1 ? lvtReg_289 : _GEN_5408; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5410 = 10'h122 == io_rdAddr_1 ? lvtReg_290 : _GEN_5409; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5411 = 10'h123 == io_rdAddr_1 ? lvtReg_291 : _GEN_5410; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5412 = 10'h124 == io_rdAddr_1 ? lvtReg_292 : _GEN_5411; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5413 = 10'h125 == io_rdAddr_1 ? lvtReg_293 : _GEN_5412; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5414 = 10'h126 == io_rdAddr_1 ? lvtReg_294 : _GEN_5413; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5415 = 10'h127 == io_rdAddr_1 ? lvtReg_295 : _GEN_5414; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5416 = 10'h128 == io_rdAddr_1 ? lvtReg_296 : _GEN_5415; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5417 = 10'h129 == io_rdAddr_1 ? lvtReg_297 : _GEN_5416; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5418 = 10'h12a == io_rdAddr_1 ? lvtReg_298 : _GEN_5417; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5419 = 10'h12b == io_rdAddr_1 ? lvtReg_299 : _GEN_5418; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5420 = 10'h12c == io_rdAddr_1 ? lvtReg_300 : _GEN_5419; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5421 = 10'h12d == io_rdAddr_1 ? lvtReg_301 : _GEN_5420; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5422 = 10'h12e == io_rdAddr_1 ? lvtReg_302 : _GEN_5421; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5423 = 10'h12f == io_rdAddr_1 ? lvtReg_303 : _GEN_5422; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5424 = 10'h130 == io_rdAddr_1 ? lvtReg_304 : _GEN_5423; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5425 = 10'h131 == io_rdAddr_1 ? lvtReg_305 : _GEN_5424; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5426 = 10'h132 == io_rdAddr_1 ? lvtReg_306 : _GEN_5425; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5427 = 10'h133 == io_rdAddr_1 ? lvtReg_307 : _GEN_5426; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5428 = 10'h134 == io_rdAddr_1 ? lvtReg_308 : _GEN_5427; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5429 = 10'h135 == io_rdAddr_1 ? lvtReg_309 : _GEN_5428; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5430 = 10'h136 == io_rdAddr_1 ? lvtReg_310 : _GEN_5429; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5431 = 10'h137 == io_rdAddr_1 ? lvtReg_311 : _GEN_5430; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5432 = 10'h138 == io_rdAddr_1 ? lvtReg_312 : _GEN_5431; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5433 = 10'h139 == io_rdAddr_1 ? lvtReg_313 : _GEN_5432; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5434 = 10'h13a == io_rdAddr_1 ? lvtReg_314 : _GEN_5433; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5435 = 10'h13b == io_rdAddr_1 ? lvtReg_315 : _GEN_5434; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5436 = 10'h13c == io_rdAddr_1 ? lvtReg_316 : _GEN_5435; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5437 = 10'h13d == io_rdAddr_1 ? lvtReg_317 : _GEN_5436; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5438 = 10'h13e == io_rdAddr_1 ? lvtReg_318 : _GEN_5437; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5439 = 10'h13f == io_rdAddr_1 ? lvtReg_319 : _GEN_5438; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5440 = 10'h140 == io_rdAddr_1 ? lvtReg_320 : _GEN_5439; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5441 = 10'h141 == io_rdAddr_1 ? lvtReg_321 : _GEN_5440; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5442 = 10'h142 == io_rdAddr_1 ? lvtReg_322 : _GEN_5441; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5443 = 10'h143 == io_rdAddr_1 ? lvtReg_323 : _GEN_5442; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5444 = 10'h144 == io_rdAddr_1 ? lvtReg_324 : _GEN_5443; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5445 = 10'h145 == io_rdAddr_1 ? lvtReg_325 : _GEN_5444; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5446 = 10'h146 == io_rdAddr_1 ? lvtReg_326 : _GEN_5445; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5447 = 10'h147 == io_rdAddr_1 ? lvtReg_327 : _GEN_5446; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5448 = 10'h148 == io_rdAddr_1 ? lvtReg_328 : _GEN_5447; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5449 = 10'h149 == io_rdAddr_1 ? lvtReg_329 : _GEN_5448; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5450 = 10'h14a == io_rdAddr_1 ? lvtReg_330 : _GEN_5449; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5451 = 10'h14b == io_rdAddr_1 ? lvtReg_331 : _GEN_5450; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5452 = 10'h14c == io_rdAddr_1 ? lvtReg_332 : _GEN_5451; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5453 = 10'h14d == io_rdAddr_1 ? lvtReg_333 : _GEN_5452; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5454 = 10'h14e == io_rdAddr_1 ? lvtReg_334 : _GEN_5453; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5455 = 10'h14f == io_rdAddr_1 ? lvtReg_335 : _GEN_5454; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5456 = 10'h150 == io_rdAddr_1 ? lvtReg_336 : _GEN_5455; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5457 = 10'h151 == io_rdAddr_1 ? lvtReg_337 : _GEN_5456; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5458 = 10'h152 == io_rdAddr_1 ? lvtReg_338 : _GEN_5457; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5459 = 10'h153 == io_rdAddr_1 ? lvtReg_339 : _GEN_5458; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5460 = 10'h154 == io_rdAddr_1 ? lvtReg_340 : _GEN_5459; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5461 = 10'h155 == io_rdAddr_1 ? lvtReg_341 : _GEN_5460; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5462 = 10'h156 == io_rdAddr_1 ? lvtReg_342 : _GEN_5461; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5463 = 10'h157 == io_rdAddr_1 ? lvtReg_343 : _GEN_5462; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5464 = 10'h158 == io_rdAddr_1 ? lvtReg_344 : _GEN_5463; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5465 = 10'h159 == io_rdAddr_1 ? lvtReg_345 : _GEN_5464; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5466 = 10'h15a == io_rdAddr_1 ? lvtReg_346 : _GEN_5465; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5467 = 10'h15b == io_rdAddr_1 ? lvtReg_347 : _GEN_5466; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5468 = 10'h15c == io_rdAddr_1 ? lvtReg_348 : _GEN_5467; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5469 = 10'h15d == io_rdAddr_1 ? lvtReg_349 : _GEN_5468; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5470 = 10'h15e == io_rdAddr_1 ? lvtReg_350 : _GEN_5469; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5471 = 10'h15f == io_rdAddr_1 ? lvtReg_351 : _GEN_5470; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5472 = 10'h160 == io_rdAddr_1 ? lvtReg_352 : _GEN_5471; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5473 = 10'h161 == io_rdAddr_1 ? lvtReg_353 : _GEN_5472; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5474 = 10'h162 == io_rdAddr_1 ? lvtReg_354 : _GEN_5473; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5475 = 10'h163 == io_rdAddr_1 ? lvtReg_355 : _GEN_5474; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5476 = 10'h164 == io_rdAddr_1 ? lvtReg_356 : _GEN_5475; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5477 = 10'h165 == io_rdAddr_1 ? lvtReg_357 : _GEN_5476; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5478 = 10'h166 == io_rdAddr_1 ? lvtReg_358 : _GEN_5477; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5479 = 10'h167 == io_rdAddr_1 ? lvtReg_359 : _GEN_5478; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5480 = 10'h168 == io_rdAddr_1 ? lvtReg_360 : _GEN_5479; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5481 = 10'h169 == io_rdAddr_1 ? lvtReg_361 : _GEN_5480; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5482 = 10'h16a == io_rdAddr_1 ? lvtReg_362 : _GEN_5481; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5483 = 10'h16b == io_rdAddr_1 ? lvtReg_363 : _GEN_5482; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5484 = 10'h16c == io_rdAddr_1 ? lvtReg_364 : _GEN_5483; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5485 = 10'h16d == io_rdAddr_1 ? lvtReg_365 : _GEN_5484; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5486 = 10'h16e == io_rdAddr_1 ? lvtReg_366 : _GEN_5485; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5487 = 10'h16f == io_rdAddr_1 ? lvtReg_367 : _GEN_5486; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5488 = 10'h170 == io_rdAddr_1 ? lvtReg_368 : _GEN_5487; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5489 = 10'h171 == io_rdAddr_1 ? lvtReg_369 : _GEN_5488; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5490 = 10'h172 == io_rdAddr_1 ? lvtReg_370 : _GEN_5489; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5491 = 10'h173 == io_rdAddr_1 ? lvtReg_371 : _GEN_5490; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5492 = 10'h174 == io_rdAddr_1 ? lvtReg_372 : _GEN_5491; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5493 = 10'h175 == io_rdAddr_1 ? lvtReg_373 : _GEN_5492; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5494 = 10'h176 == io_rdAddr_1 ? lvtReg_374 : _GEN_5493; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5495 = 10'h177 == io_rdAddr_1 ? lvtReg_375 : _GEN_5494; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5496 = 10'h178 == io_rdAddr_1 ? lvtReg_376 : _GEN_5495; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5497 = 10'h179 == io_rdAddr_1 ? lvtReg_377 : _GEN_5496; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5498 = 10'h17a == io_rdAddr_1 ? lvtReg_378 : _GEN_5497; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5499 = 10'h17b == io_rdAddr_1 ? lvtReg_379 : _GEN_5498; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5500 = 10'h17c == io_rdAddr_1 ? lvtReg_380 : _GEN_5499; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5501 = 10'h17d == io_rdAddr_1 ? lvtReg_381 : _GEN_5500; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5502 = 10'h17e == io_rdAddr_1 ? lvtReg_382 : _GEN_5501; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5503 = 10'h17f == io_rdAddr_1 ? lvtReg_383 : _GEN_5502; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5504 = 10'h180 == io_rdAddr_1 ? lvtReg_384 : _GEN_5503; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5505 = 10'h181 == io_rdAddr_1 ? lvtReg_385 : _GEN_5504; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5506 = 10'h182 == io_rdAddr_1 ? lvtReg_386 : _GEN_5505; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5507 = 10'h183 == io_rdAddr_1 ? lvtReg_387 : _GEN_5506; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5508 = 10'h184 == io_rdAddr_1 ? lvtReg_388 : _GEN_5507; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5509 = 10'h185 == io_rdAddr_1 ? lvtReg_389 : _GEN_5508; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5510 = 10'h186 == io_rdAddr_1 ? lvtReg_390 : _GEN_5509; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5511 = 10'h187 == io_rdAddr_1 ? lvtReg_391 : _GEN_5510; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5512 = 10'h188 == io_rdAddr_1 ? lvtReg_392 : _GEN_5511; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5513 = 10'h189 == io_rdAddr_1 ? lvtReg_393 : _GEN_5512; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5514 = 10'h18a == io_rdAddr_1 ? lvtReg_394 : _GEN_5513; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5515 = 10'h18b == io_rdAddr_1 ? lvtReg_395 : _GEN_5514; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5516 = 10'h18c == io_rdAddr_1 ? lvtReg_396 : _GEN_5515; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5517 = 10'h18d == io_rdAddr_1 ? lvtReg_397 : _GEN_5516; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5518 = 10'h18e == io_rdAddr_1 ? lvtReg_398 : _GEN_5517; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5519 = 10'h18f == io_rdAddr_1 ? lvtReg_399 : _GEN_5518; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5520 = 10'h190 == io_rdAddr_1 ? lvtReg_400 : _GEN_5519; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5521 = 10'h191 == io_rdAddr_1 ? lvtReg_401 : _GEN_5520; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5522 = 10'h192 == io_rdAddr_1 ? lvtReg_402 : _GEN_5521; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5523 = 10'h193 == io_rdAddr_1 ? lvtReg_403 : _GEN_5522; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5524 = 10'h194 == io_rdAddr_1 ? lvtReg_404 : _GEN_5523; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5525 = 10'h195 == io_rdAddr_1 ? lvtReg_405 : _GEN_5524; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5526 = 10'h196 == io_rdAddr_1 ? lvtReg_406 : _GEN_5525; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5527 = 10'h197 == io_rdAddr_1 ? lvtReg_407 : _GEN_5526; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5528 = 10'h198 == io_rdAddr_1 ? lvtReg_408 : _GEN_5527; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5529 = 10'h199 == io_rdAddr_1 ? lvtReg_409 : _GEN_5528; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5530 = 10'h19a == io_rdAddr_1 ? lvtReg_410 : _GEN_5529; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5531 = 10'h19b == io_rdAddr_1 ? lvtReg_411 : _GEN_5530; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5532 = 10'h19c == io_rdAddr_1 ? lvtReg_412 : _GEN_5531; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5533 = 10'h19d == io_rdAddr_1 ? lvtReg_413 : _GEN_5532; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5534 = 10'h19e == io_rdAddr_1 ? lvtReg_414 : _GEN_5533; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5535 = 10'h19f == io_rdAddr_1 ? lvtReg_415 : _GEN_5534; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5536 = 10'h1a0 == io_rdAddr_1 ? lvtReg_416 : _GEN_5535; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5537 = 10'h1a1 == io_rdAddr_1 ? lvtReg_417 : _GEN_5536; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5538 = 10'h1a2 == io_rdAddr_1 ? lvtReg_418 : _GEN_5537; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5539 = 10'h1a3 == io_rdAddr_1 ? lvtReg_419 : _GEN_5538; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5540 = 10'h1a4 == io_rdAddr_1 ? lvtReg_420 : _GEN_5539; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5541 = 10'h1a5 == io_rdAddr_1 ? lvtReg_421 : _GEN_5540; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5542 = 10'h1a6 == io_rdAddr_1 ? lvtReg_422 : _GEN_5541; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5543 = 10'h1a7 == io_rdAddr_1 ? lvtReg_423 : _GEN_5542; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5544 = 10'h1a8 == io_rdAddr_1 ? lvtReg_424 : _GEN_5543; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5545 = 10'h1a9 == io_rdAddr_1 ? lvtReg_425 : _GEN_5544; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5546 = 10'h1aa == io_rdAddr_1 ? lvtReg_426 : _GEN_5545; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5547 = 10'h1ab == io_rdAddr_1 ? lvtReg_427 : _GEN_5546; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5548 = 10'h1ac == io_rdAddr_1 ? lvtReg_428 : _GEN_5547; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5549 = 10'h1ad == io_rdAddr_1 ? lvtReg_429 : _GEN_5548; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5550 = 10'h1ae == io_rdAddr_1 ? lvtReg_430 : _GEN_5549; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5551 = 10'h1af == io_rdAddr_1 ? lvtReg_431 : _GEN_5550; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5552 = 10'h1b0 == io_rdAddr_1 ? lvtReg_432 : _GEN_5551; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5553 = 10'h1b1 == io_rdAddr_1 ? lvtReg_433 : _GEN_5552; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5554 = 10'h1b2 == io_rdAddr_1 ? lvtReg_434 : _GEN_5553; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5555 = 10'h1b3 == io_rdAddr_1 ? lvtReg_435 : _GEN_5554; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5556 = 10'h1b4 == io_rdAddr_1 ? lvtReg_436 : _GEN_5555; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5557 = 10'h1b5 == io_rdAddr_1 ? lvtReg_437 : _GEN_5556; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5558 = 10'h1b6 == io_rdAddr_1 ? lvtReg_438 : _GEN_5557; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5559 = 10'h1b7 == io_rdAddr_1 ? lvtReg_439 : _GEN_5558; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5560 = 10'h1b8 == io_rdAddr_1 ? lvtReg_440 : _GEN_5559; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5561 = 10'h1b9 == io_rdAddr_1 ? lvtReg_441 : _GEN_5560; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5562 = 10'h1ba == io_rdAddr_1 ? lvtReg_442 : _GEN_5561; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5563 = 10'h1bb == io_rdAddr_1 ? lvtReg_443 : _GEN_5562; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5564 = 10'h1bc == io_rdAddr_1 ? lvtReg_444 : _GEN_5563; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5565 = 10'h1bd == io_rdAddr_1 ? lvtReg_445 : _GEN_5564; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5566 = 10'h1be == io_rdAddr_1 ? lvtReg_446 : _GEN_5565; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5567 = 10'h1bf == io_rdAddr_1 ? lvtReg_447 : _GEN_5566; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5568 = 10'h1c0 == io_rdAddr_1 ? lvtReg_448 : _GEN_5567; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5569 = 10'h1c1 == io_rdAddr_1 ? lvtReg_449 : _GEN_5568; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5570 = 10'h1c2 == io_rdAddr_1 ? lvtReg_450 : _GEN_5569; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5571 = 10'h1c3 == io_rdAddr_1 ? lvtReg_451 : _GEN_5570; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5572 = 10'h1c4 == io_rdAddr_1 ? lvtReg_452 : _GEN_5571; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5573 = 10'h1c5 == io_rdAddr_1 ? lvtReg_453 : _GEN_5572; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5574 = 10'h1c6 == io_rdAddr_1 ? lvtReg_454 : _GEN_5573; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5575 = 10'h1c7 == io_rdAddr_1 ? lvtReg_455 : _GEN_5574; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5576 = 10'h1c8 == io_rdAddr_1 ? lvtReg_456 : _GEN_5575; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5577 = 10'h1c9 == io_rdAddr_1 ? lvtReg_457 : _GEN_5576; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5578 = 10'h1ca == io_rdAddr_1 ? lvtReg_458 : _GEN_5577; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5579 = 10'h1cb == io_rdAddr_1 ? lvtReg_459 : _GEN_5578; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5580 = 10'h1cc == io_rdAddr_1 ? lvtReg_460 : _GEN_5579; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5581 = 10'h1cd == io_rdAddr_1 ? lvtReg_461 : _GEN_5580; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5582 = 10'h1ce == io_rdAddr_1 ? lvtReg_462 : _GEN_5581; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5583 = 10'h1cf == io_rdAddr_1 ? lvtReg_463 : _GEN_5582; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5584 = 10'h1d0 == io_rdAddr_1 ? lvtReg_464 : _GEN_5583; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5585 = 10'h1d1 == io_rdAddr_1 ? lvtReg_465 : _GEN_5584; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5586 = 10'h1d2 == io_rdAddr_1 ? lvtReg_466 : _GEN_5585; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5587 = 10'h1d3 == io_rdAddr_1 ? lvtReg_467 : _GEN_5586; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5588 = 10'h1d4 == io_rdAddr_1 ? lvtReg_468 : _GEN_5587; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5589 = 10'h1d5 == io_rdAddr_1 ? lvtReg_469 : _GEN_5588; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5590 = 10'h1d6 == io_rdAddr_1 ? lvtReg_470 : _GEN_5589; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5591 = 10'h1d7 == io_rdAddr_1 ? lvtReg_471 : _GEN_5590; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5592 = 10'h1d8 == io_rdAddr_1 ? lvtReg_472 : _GEN_5591; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5593 = 10'h1d9 == io_rdAddr_1 ? lvtReg_473 : _GEN_5592; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5594 = 10'h1da == io_rdAddr_1 ? lvtReg_474 : _GEN_5593; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5595 = 10'h1db == io_rdAddr_1 ? lvtReg_475 : _GEN_5594; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5596 = 10'h1dc == io_rdAddr_1 ? lvtReg_476 : _GEN_5595; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5597 = 10'h1dd == io_rdAddr_1 ? lvtReg_477 : _GEN_5596; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5598 = 10'h1de == io_rdAddr_1 ? lvtReg_478 : _GEN_5597; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5599 = 10'h1df == io_rdAddr_1 ? lvtReg_479 : _GEN_5598; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5600 = 10'h1e0 == io_rdAddr_1 ? lvtReg_480 : _GEN_5599; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5601 = 10'h1e1 == io_rdAddr_1 ? lvtReg_481 : _GEN_5600; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5602 = 10'h1e2 == io_rdAddr_1 ? lvtReg_482 : _GEN_5601; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5603 = 10'h1e3 == io_rdAddr_1 ? lvtReg_483 : _GEN_5602; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5604 = 10'h1e4 == io_rdAddr_1 ? lvtReg_484 : _GEN_5603; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5605 = 10'h1e5 == io_rdAddr_1 ? lvtReg_485 : _GEN_5604; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5606 = 10'h1e6 == io_rdAddr_1 ? lvtReg_486 : _GEN_5605; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5607 = 10'h1e7 == io_rdAddr_1 ? lvtReg_487 : _GEN_5606; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5608 = 10'h1e8 == io_rdAddr_1 ? lvtReg_488 : _GEN_5607; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5609 = 10'h1e9 == io_rdAddr_1 ? lvtReg_489 : _GEN_5608; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5610 = 10'h1ea == io_rdAddr_1 ? lvtReg_490 : _GEN_5609; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5611 = 10'h1eb == io_rdAddr_1 ? lvtReg_491 : _GEN_5610; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5612 = 10'h1ec == io_rdAddr_1 ? lvtReg_492 : _GEN_5611; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5613 = 10'h1ed == io_rdAddr_1 ? lvtReg_493 : _GEN_5612; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5614 = 10'h1ee == io_rdAddr_1 ? lvtReg_494 : _GEN_5613; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5615 = 10'h1ef == io_rdAddr_1 ? lvtReg_495 : _GEN_5614; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5616 = 10'h1f0 == io_rdAddr_1 ? lvtReg_496 : _GEN_5615; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5617 = 10'h1f1 == io_rdAddr_1 ? lvtReg_497 : _GEN_5616; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5618 = 10'h1f2 == io_rdAddr_1 ? lvtReg_498 : _GEN_5617; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5619 = 10'h1f3 == io_rdAddr_1 ? lvtReg_499 : _GEN_5618; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5620 = 10'h1f4 == io_rdAddr_1 ? lvtReg_500 : _GEN_5619; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5621 = 10'h1f5 == io_rdAddr_1 ? lvtReg_501 : _GEN_5620; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5622 = 10'h1f6 == io_rdAddr_1 ? lvtReg_502 : _GEN_5621; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5623 = 10'h1f7 == io_rdAddr_1 ? lvtReg_503 : _GEN_5622; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5624 = 10'h1f8 == io_rdAddr_1 ? lvtReg_504 : _GEN_5623; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5625 = 10'h1f9 == io_rdAddr_1 ? lvtReg_505 : _GEN_5624; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5626 = 10'h1fa == io_rdAddr_1 ? lvtReg_506 : _GEN_5625; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5627 = 10'h1fb == io_rdAddr_1 ? lvtReg_507 : _GEN_5626; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5628 = 10'h1fc == io_rdAddr_1 ? lvtReg_508 : _GEN_5627; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5629 = 10'h1fd == io_rdAddr_1 ? lvtReg_509 : _GEN_5628; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5630 = 10'h1fe == io_rdAddr_1 ? lvtReg_510 : _GEN_5629; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5631 = 10'h1ff == io_rdAddr_1 ? lvtReg_511 : _GEN_5630; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5632 = 10'h200 == io_rdAddr_1 ? lvtReg_512 : _GEN_5631; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5633 = 10'h201 == io_rdAddr_1 ? lvtReg_513 : _GEN_5632; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5634 = 10'h202 == io_rdAddr_1 ? lvtReg_514 : _GEN_5633; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5635 = 10'h203 == io_rdAddr_1 ? lvtReg_515 : _GEN_5634; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5636 = 10'h204 == io_rdAddr_1 ? lvtReg_516 : _GEN_5635; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5637 = 10'h205 == io_rdAddr_1 ? lvtReg_517 : _GEN_5636; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5638 = 10'h206 == io_rdAddr_1 ? lvtReg_518 : _GEN_5637; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5639 = 10'h207 == io_rdAddr_1 ? lvtReg_519 : _GEN_5638; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5640 = 10'h208 == io_rdAddr_1 ? lvtReg_520 : _GEN_5639; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5641 = 10'h209 == io_rdAddr_1 ? lvtReg_521 : _GEN_5640; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5642 = 10'h20a == io_rdAddr_1 ? lvtReg_522 : _GEN_5641; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5643 = 10'h20b == io_rdAddr_1 ? lvtReg_523 : _GEN_5642; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5644 = 10'h20c == io_rdAddr_1 ? lvtReg_524 : _GEN_5643; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5645 = 10'h20d == io_rdAddr_1 ? lvtReg_525 : _GEN_5644; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5646 = 10'h20e == io_rdAddr_1 ? lvtReg_526 : _GEN_5645; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5647 = 10'h20f == io_rdAddr_1 ? lvtReg_527 : _GEN_5646; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5648 = 10'h210 == io_rdAddr_1 ? lvtReg_528 : _GEN_5647; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5649 = 10'h211 == io_rdAddr_1 ? lvtReg_529 : _GEN_5648; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5650 = 10'h212 == io_rdAddr_1 ? lvtReg_530 : _GEN_5649; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5651 = 10'h213 == io_rdAddr_1 ? lvtReg_531 : _GEN_5650; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5652 = 10'h214 == io_rdAddr_1 ? lvtReg_532 : _GEN_5651; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5653 = 10'h215 == io_rdAddr_1 ? lvtReg_533 : _GEN_5652; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5654 = 10'h216 == io_rdAddr_1 ? lvtReg_534 : _GEN_5653; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5655 = 10'h217 == io_rdAddr_1 ? lvtReg_535 : _GEN_5654; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5656 = 10'h218 == io_rdAddr_1 ? lvtReg_536 : _GEN_5655; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5657 = 10'h219 == io_rdAddr_1 ? lvtReg_537 : _GEN_5656; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5658 = 10'h21a == io_rdAddr_1 ? lvtReg_538 : _GEN_5657; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5659 = 10'h21b == io_rdAddr_1 ? lvtReg_539 : _GEN_5658; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5660 = 10'h21c == io_rdAddr_1 ? lvtReg_540 : _GEN_5659; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5661 = 10'h21d == io_rdAddr_1 ? lvtReg_541 : _GEN_5660; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5662 = 10'h21e == io_rdAddr_1 ? lvtReg_542 : _GEN_5661; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5663 = 10'h21f == io_rdAddr_1 ? lvtReg_543 : _GEN_5662; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5664 = 10'h220 == io_rdAddr_1 ? lvtReg_544 : _GEN_5663; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5665 = 10'h221 == io_rdAddr_1 ? lvtReg_545 : _GEN_5664; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5666 = 10'h222 == io_rdAddr_1 ? lvtReg_546 : _GEN_5665; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5667 = 10'h223 == io_rdAddr_1 ? lvtReg_547 : _GEN_5666; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5668 = 10'h224 == io_rdAddr_1 ? lvtReg_548 : _GEN_5667; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5669 = 10'h225 == io_rdAddr_1 ? lvtReg_549 : _GEN_5668; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5670 = 10'h226 == io_rdAddr_1 ? lvtReg_550 : _GEN_5669; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5671 = 10'h227 == io_rdAddr_1 ? lvtReg_551 : _GEN_5670; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5672 = 10'h228 == io_rdAddr_1 ? lvtReg_552 : _GEN_5671; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5673 = 10'h229 == io_rdAddr_1 ? lvtReg_553 : _GEN_5672; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5674 = 10'h22a == io_rdAddr_1 ? lvtReg_554 : _GEN_5673; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5675 = 10'h22b == io_rdAddr_1 ? lvtReg_555 : _GEN_5674; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5676 = 10'h22c == io_rdAddr_1 ? lvtReg_556 : _GEN_5675; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5677 = 10'h22d == io_rdAddr_1 ? lvtReg_557 : _GEN_5676; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5678 = 10'h22e == io_rdAddr_1 ? lvtReg_558 : _GEN_5677; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5679 = 10'h22f == io_rdAddr_1 ? lvtReg_559 : _GEN_5678; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5680 = 10'h230 == io_rdAddr_1 ? lvtReg_560 : _GEN_5679; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5681 = 10'h231 == io_rdAddr_1 ? lvtReg_561 : _GEN_5680; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5682 = 10'h232 == io_rdAddr_1 ? lvtReg_562 : _GEN_5681; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5683 = 10'h233 == io_rdAddr_1 ? lvtReg_563 : _GEN_5682; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5684 = 10'h234 == io_rdAddr_1 ? lvtReg_564 : _GEN_5683; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5685 = 10'h235 == io_rdAddr_1 ? lvtReg_565 : _GEN_5684; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5686 = 10'h236 == io_rdAddr_1 ? lvtReg_566 : _GEN_5685; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5687 = 10'h237 == io_rdAddr_1 ? lvtReg_567 : _GEN_5686; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5688 = 10'h238 == io_rdAddr_1 ? lvtReg_568 : _GEN_5687; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5689 = 10'h239 == io_rdAddr_1 ? lvtReg_569 : _GEN_5688; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5690 = 10'h23a == io_rdAddr_1 ? lvtReg_570 : _GEN_5689; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5691 = 10'h23b == io_rdAddr_1 ? lvtReg_571 : _GEN_5690; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5692 = 10'h23c == io_rdAddr_1 ? lvtReg_572 : _GEN_5691; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5693 = 10'h23d == io_rdAddr_1 ? lvtReg_573 : _GEN_5692; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5694 = 10'h23e == io_rdAddr_1 ? lvtReg_574 : _GEN_5693; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5695 = 10'h23f == io_rdAddr_1 ? lvtReg_575 : _GEN_5694; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5696 = 10'h240 == io_rdAddr_1 ? lvtReg_576 : _GEN_5695; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5697 = 10'h241 == io_rdAddr_1 ? lvtReg_577 : _GEN_5696; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5698 = 10'h242 == io_rdAddr_1 ? lvtReg_578 : _GEN_5697; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5699 = 10'h243 == io_rdAddr_1 ? lvtReg_579 : _GEN_5698; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5700 = 10'h244 == io_rdAddr_1 ? lvtReg_580 : _GEN_5699; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5701 = 10'h245 == io_rdAddr_1 ? lvtReg_581 : _GEN_5700; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5702 = 10'h246 == io_rdAddr_1 ? lvtReg_582 : _GEN_5701; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5703 = 10'h247 == io_rdAddr_1 ? lvtReg_583 : _GEN_5702; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5704 = 10'h248 == io_rdAddr_1 ? lvtReg_584 : _GEN_5703; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5705 = 10'h249 == io_rdAddr_1 ? lvtReg_585 : _GEN_5704; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5706 = 10'h24a == io_rdAddr_1 ? lvtReg_586 : _GEN_5705; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5707 = 10'h24b == io_rdAddr_1 ? lvtReg_587 : _GEN_5706; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5708 = 10'h24c == io_rdAddr_1 ? lvtReg_588 : _GEN_5707; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5709 = 10'h24d == io_rdAddr_1 ? lvtReg_589 : _GEN_5708; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5710 = 10'h24e == io_rdAddr_1 ? lvtReg_590 : _GEN_5709; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5711 = 10'h24f == io_rdAddr_1 ? lvtReg_591 : _GEN_5710; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5712 = 10'h250 == io_rdAddr_1 ? lvtReg_592 : _GEN_5711; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5713 = 10'h251 == io_rdAddr_1 ? lvtReg_593 : _GEN_5712; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5714 = 10'h252 == io_rdAddr_1 ? lvtReg_594 : _GEN_5713; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5715 = 10'h253 == io_rdAddr_1 ? lvtReg_595 : _GEN_5714; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5716 = 10'h254 == io_rdAddr_1 ? lvtReg_596 : _GEN_5715; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5717 = 10'h255 == io_rdAddr_1 ? lvtReg_597 : _GEN_5716; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5718 = 10'h256 == io_rdAddr_1 ? lvtReg_598 : _GEN_5717; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5719 = 10'h257 == io_rdAddr_1 ? lvtReg_599 : _GEN_5718; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5720 = 10'h258 == io_rdAddr_1 ? lvtReg_600 : _GEN_5719; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5721 = 10'h259 == io_rdAddr_1 ? lvtReg_601 : _GEN_5720; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5722 = 10'h25a == io_rdAddr_1 ? lvtReg_602 : _GEN_5721; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5723 = 10'h25b == io_rdAddr_1 ? lvtReg_603 : _GEN_5722; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5724 = 10'h25c == io_rdAddr_1 ? lvtReg_604 : _GEN_5723; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5725 = 10'h25d == io_rdAddr_1 ? lvtReg_605 : _GEN_5724; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5726 = 10'h25e == io_rdAddr_1 ? lvtReg_606 : _GEN_5725; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5727 = 10'h25f == io_rdAddr_1 ? lvtReg_607 : _GEN_5726; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5728 = 10'h260 == io_rdAddr_1 ? lvtReg_608 : _GEN_5727; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5729 = 10'h261 == io_rdAddr_1 ? lvtReg_609 : _GEN_5728; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5730 = 10'h262 == io_rdAddr_1 ? lvtReg_610 : _GEN_5729; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5731 = 10'h263 == io_rdAddr_1 ? lvtReg_611 : _GEN_5730; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5732 = 10'h264 == io_rdAddr_1 ? lvtReg_612 : _GEN_5731; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5733 = 10'h265 == io_rdAddr_1 ? lvtReg_613 : _GEN_5732; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5734 = 10'h266 == io_rdAddr_1 ? lvtReg_614 : _GEN_5733; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5735 = 10'h267 == io_rdAddr_1 ? lvtReg_615 : _GEN_5734; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5736 = 10'h268 == io_rdAddr_1 ? lvtReg_616 : _GEN_5735; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5737 = 10'h269 == io_rdAddr_1 ? lvtReg_617 : _GEN_5736; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5738 = 10'h26a == io_rdAddr_1 ? lvtReg_618 : _GEN_5737; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5739 = 10'h26b == io_rdAddr_1 ? lvtReg_619 : _GEN_5738; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5740 = 10'h26c == io_rdAddr_1 ? lvtReg_620 : _GEN_5739; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5741 = 10'h26d == io_rdAddr_1 ? lvtReg_621 : _GEN_5740; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5742 = 10'h26e == io_rdAddr_1 ? lvtReg_622 : _GEN_5741; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5743 = 10'h26f == io_rdAddr_1 ? lvtReg_623 : _GEN_5742; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5744 = 10'h270 == io_rdAddr_1 ? lvtReg_624 : _GEN_5743; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5745 = 10'h271 == io_rdAddr_1 ? lvtReg_625 : _GEN_5744; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5746 = 10'h272 == io_rdAddr_1 ? lvtReg_626 : _GEN_5745; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5747 = 10'h273 == io_rdAddr_1 ? lvtReg_627 : _GEN_5746; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5748 = 10'h274 == io_rdAddr_1 ? lvtReg_628 : _GEN_5747; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5749 = 10'h275 == io_rdAddr_1 ? lvtReg_629 : _GEN_5748; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5750 = 10'h276 == io_rdAddr_1 ? lvtReg_630 : _GEN_5749; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5751 = 10'h277 == io_rdAddr_1 ? lvtReg_631 : _GEN_5750; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5752 = 10'h278 == io_rdAddr_1 ? lvtReg_632 : _GEN_5751; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5753 = 10'h279 == io_rdAddr_1 ? lvtReg_633 : _GEN_5752; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5754 = 10'h27a == io_rdAddr_1 ? lvtReg_634 : _GEN_5753; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5755 = 10'h27b == io_rdAddr_1 ? lvtReg_635 : _GEN_5754; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5756 = 10'h27c == io_rdAddr_1 ? lvtReg_636 : _GEN_5755; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5757 = 10'h27d == io_rdAddr_1 ? lvtReg_637 : _GEN_5756; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5758 = 10'h27e == io_rdAddr_1 ? lvtReg_638 : _GEN_5757; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5759 = 10'h27f == io_rdAddr_1 ? lvtReg_639 : _GEN_5758; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5760 = 10'h280 == io_rdAddr_1 ? lvtReg_640 : _GEN_5759; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5761 = 10'h281 == io_rdAddr_1 ? lvtReg_641 : _GEN_5760; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5762 = 10'h282 == io_rdAddr_1 ? lvtReg_642 : _GEN_5761; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5763 = 10'h283 == io_rdAddr_1 ? lvtReg_643 : _GEN_5762; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5764 = 10'h284 == io_rdAddr_1 ? lvtReg_644 : _GEN_5763; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5765 = 10'h285 == io_rdAddr_1 ? lvtReg_645 : _GEN_5764; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5766 = 10'h286 == io_rdAddr_1 ? lvtReg_646 : _GEN_5765; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5767 = 10'h287 == io_rdAddr_1 ? lvtReg_647 : _GEN_5766; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5768 = 10'h288 == io_rdAddr_1 ? lvtReg_648 : _GEN_5767; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5769 = 10'h289 == io_rdAddr_1 ? lvtReg_649 : _GEN_5768; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5770 = 10'h28a == io_rdAddr_1 ? lvtReg_650 : _GEN_5769; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5771 = 10'h28b == io_rdAddr_1 ? lvtReg_651 : _GEN_5770; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5772 = 10'h28c == io_rdAddr_1 ? lvtReg_652 : _GEN_5771; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5773 = 10'h28d == io_rdAddr_1 ? lvtReg_653 : _GEN_5772; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5774 = 10'h28e == io_rdAddr_1 ? lvtReg_654 : _GEN_5773; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5775 = 10'h28f == io_rdAddr_1 ? lvtReg_655 : _GEN_5774; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5776 = 10'h290 == io_rdAddr_1 ? lvtReg_656 : _GEN_5775; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5777 = 10'h291 == io_rdAddr_1 ? lvtReg_657 : _GEN_5776; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5778 = 10'h292 == io_rdAddr_1 ? lvtReg_658 : _GEN_5777; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5779 = 10'h293 == io_rdAddr_1 ? lvtReg_659 : _GEN_5778; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5780 = 10'h294 == io_rdAddr_1 ? lvtReg_660 : _GEN_5779; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5781 = 10'h295 == io_rdAddr_1 ? lvtReg_661 : _GEN_5780; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5782 = 10'h296 == io_rdAddr_1 ? lvtReg_662 : _GEN_5781; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5783 = 10'h297 == io_rdAddr_1 ? lvtReg_663 : _GEN_5782; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5784 = 10'h298 == io_rdAddr_1 ? lvtReg_664 : _GEN_5783; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5785 = 10'h299 == io_rdAddr_1 ? lvtReg_665 : _GEN_5784; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5786 = 10'h29a == io_rdAddr_1 ? lvtReg_666 : _GEN_5785; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5787 = 10'h29b == io_rdAddr_1 ? lvtReg_667 : _GEN_5786; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5788 = 10'h29c == io_rdAddr_1 ? lvtReg_668 : _GEN_5787; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5789 = 10'h29d == io_rdAddr_1 ? lvtReg_669 : _GEN_5788; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5790 = 10'h29e == io_rdAddr_1 ? lvtReg_670 : _GEN_5789; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5791 = 10'h29f == io_rdAddr_1 ? lvtReg_671 : _GEN_5790; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5792 = 10'h2a0 == io_rdAddr_1 ? lvtReg_672 : _GEN_5791; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5793 = 10'h2a1 == io_rdAddr_1 ? lvtReg_673 : _GEN_5792; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5794 = 10'h2a2 == io_rdAddr_1 ? lvtReg_674 : _GEN_5793; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5795 = 10'h2a3 == io_rdAddr_1 ? lvtReg_675 : _GEN_5794; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5796 = 10'h2a4 == io_rdAddr_1 ? lvtReg_676 : _GEN_5795; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5797 = 10'h2a5 == io_rdAddr_1 ? lvtReg_677 : _GEN_5796; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5798 = 10'h2a6 == io_rdAddr_1 ? lvtReg_678 : _GEN_5797; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5799 = 10'h2a7 == io_rdAddr_1 ? lvtReg_679 : _GEN_5798; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5800 = 10'h2a8 == io_rdAddr_1 ? lvtReg_680 : _GEN_5799; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5801 = 10'h2a9 == io_rdAddr_1 ? lvtReg_681 : _GEN_5800; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5802 = 10'h2aa == io_rdAddr_1 ? lvtReg_682 : _GEN_5801; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5803 = 10'h2ab == io_rdAddr_1 ? lvtReg_683 : _GEN_5802; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5804 = 10'h2ac == io_rdAddr_1 ? lvtReg_684 : _GEN_5803; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5805 = 10'h2ad == io_rdAddr_1 ? lvtReg_685 : _GEN_5804; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5806 = 10'h2ae == io_rdAddr_1 ? lvtReg_686 : _GEN_5805; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5807 = 10'h2af == io_rdAddr_1 ? lvtReg_687 : _GEN_5806; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5808 = 10'h2b0 == io_rdAddr_1 ? lvtReg_688 : _GEN_5807; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5809 = 10'h2b1 == io_rdAddr_1 ? lvtReg_689 : _GEN_5808; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5810 = 10'h2b2 == io_rdAddr_1 ? lvtReg_690 : _GEN_5809; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5811 = 10'h2b3 == io_rdAddr_1 ? lvtReg_691 : _GEN_5810; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5812 = 10'h2b4 == io_rdAddr_1 ? lvtReg_692 : _GEN_5811; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5813 = 10'h2b5 == io_rdAddr_1 ? lvtReg_693 : _GEN_5812; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5814 = 10'h2b6 == io_rdAddr_1 ? lvtReg_694 : _GEN_5813; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5815 = 10'h2b7 == io_rdAddr_1 ? lvtReg_695 : _GEN_5814; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5816 = 10'h2b8 == io_rdAddr_1 ? lvtReg_696 : _GEN_5815; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5817 = 10'h2b9 == io_rdAddr_1 ? lvtReg_697 : _GEN_5816; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5818 = 10'h2ba == io_rdAddr_1 ? lvtReg_698 : _GEN_5817; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5819 = 10'h2bb == io_rdAddr_1 ? lvtReg_699 : _GEN_5818; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5820 = 10'h2bc == io_rdAddr_1 ? lvtReg_700 : _GEN_5819; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5821 = 10'h2bd == io_rdAddr_1 ? lvtReg_701 : _GEN_5820; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5822 = 10'h2be == io_rdAddr_1 ? lvtReg_702 : _GEN_5821; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5823 = 10'h2bf == io_rdAddr_1 ? lvtReg_703 : _GEN_5822; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5824 = 10'h2c0 == io_rdAddr_1 ? lvtReg_704 : _GEN_5823; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5825 = 10'h2c1 == io_rdAddr_1 ? lvtReg_705 : _GEN_5824; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5826 = 10'h2c2 == io_rdAddr_1 ? lvtReg_706 : _GEN_5825; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5827 = 10'h2c3 == io_rdAddr_1 ? lvtReg_707 : _GEN_5826; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5828 = 10'h2c4 == io_rdAddr_1 ? lvtReg_708 : _GEN_5827; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5829 = 10'h2c5 == io_rdAddr_1 ? lvtReg_709 : _GEN_5828; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5830 = 10'h2c6 == io_rdAddr_1 ? lvtReg_710 : _GEN_5829; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5831 = 10'h2c7 == io_rdAddr_1 ? lvtReg_711 : _GEN_5830; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5832 = 10'h2c8 == io_rdAddr_1 ? lvtReg_712 : _GEN_5831; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5833 = 10'h2c9 == io_rdAddr_1 ? lvtReg_713 : _GEN_5832; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5834 = 10'h2ca == io_rdAddr_1 ? lvtReg_714 : _GEN_5833; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5835 = 10'h2cb == io_rdAddr_1 ? lvtReg_715 : _GEN_5834; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5836 = 10'h2cc == io_rdAddr_1 ? lvtReg_716 : _GEN_5835; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5837 = 10'h2cd == io_rdAddr_1 ? lvtReg_717 : _GEN_5836; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5838 = 10'h2ce == io_rdAddr_1 ? lvtReg_718 : _GEN_5837; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5839 = 10'h2cf == io_rdAddr_1 ? lvtReg_719 : _GEN_5838; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5840 = 10'h2d0 == io_rdAddr_1 ? lvtReg_720 : _GEN_5839; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5841 = 10'h2d1 == io_rdAddr_1 ? lvtReg_721 : _GEN_5840; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5842 = 10'h2d2 == io_rdAddr_1 ? lvtReg_722 : _GEN_5841; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5843 = 10'h2d3 == io_rdAddr_1 ? lvtReg_723 : _GEN_5842; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5844 = 10'h2d4 == io_rdAddr_1 ? lvtReg_724 : _GEN_5843; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5845 = 10'h2d5 == io_rdAddr_1 ? lvtReg_725 : _GEN_5844; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5846 = 10'h2d6 == io_rdAddr_1 ? lvtReg_726 : _GEN_5845; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5847 = 10'h2d7 == io_rdAddr_1 ? lvtReg_727 : _GEN_5846; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5848 = 10'h2d8 == io_rdAddr_1 ? lvtReg_728 : _GEN_5847; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5849 = 10'h2d9 == io_rdAddr_1 ? lvtReg_729 : _GEN_5848; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5850 = 10'h2da == io_rdAddr_1 ? lvtReg_730 : _GEN_5849; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5851 = 10'h2db == io_rdAddr_1 ? lvtReg_731 : _GEN_5850; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5852 = 10'h2dc == io_rdAddr_1 ? lvtReg_732 : _GEN_5851; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5853 = 10'h2dd == io_rdAddr_1 ? lvtReg_733 : _GEN_5852; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5854 = 10'h2de == io_rdAddr_1 ? lvtReg_734 : _GEN_5853; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5855 = 10'h2df == io_rdAddr_1 ? lvtReg_735 : _GEN_5854; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5856 = 10'h2e0 == io_rdAddr_1 ? lvtReg_736 : _GEN_5855; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5857 = 10'h2e1 == io_rdAddr_1 ? lvtReg_737 : _GEN_5856; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5858 = 10'h2e2 == io_rdAddr_1 ? lvtReg_738 : _GEN_5857; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5859 = 10'h2e3 == io_rdAddr_1 ? lvtReg_739 : _GEN_5858; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5860 = 10'h2e4 == io_rdAddr_1 ? lvtReg_740 : _GEN_5859; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5861 = 10'h2e5 == io_rdAddr_1 ? lvtReg_741 : _GEN_5860; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5862 = 10'h2e6 == io_rdAddr_1 ? lvtReg_742 : _GEN_5861; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5863 = 10'h2e7 == io_rdAddr_1 ? lvtReg_743 : _GEN_5862; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5864 = 10'h2e8 == io_rdAddr_1 ? lvtReg_744 : _GEN_5863; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5865 = 10'h2e9 == io_rdAddr_1 ? lvtReg_745 : _GEN_5864; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5866 = 10'h2ea == io_rdAddr_1 ? lvtReg_746 : _GEN_5865; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5867 = 10'h2eb == io_rdAddr_1 ? lvtReg_747 : _GEN_5866; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5868 = 10'h2ec == io_rdAddr_1 ? lvtReg_748 : _GEN_5867; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5869 = 10'h2ed == io_rdAddr_1 ? lvtReg_749 : _GEN_5868; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5870 = 10'h2ee == io_rdAddr_1 ? lvtReg_750 : _GEN_5869; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5871 = 10'h2ef == io_rdAddr_1 ? lvtReg_751 : _GEN_5870; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5872 = 10'h2f0 == io_rdAddr_1 ? lvtReg_752 : _GEN_5871; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5873 = 10'h2f1 == io_rdAddr_1 ? lvtReg_753 : _GEN_5872; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5874 = 10'h2f2 == io_rdAddr_1 ? lvtReg_754 : _GEN_5873; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5875 = 10'h2f3 == io_rdAddr_1 ? lvtReg_755 : _GEN_5874; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5876 = 10'h2f4 == io_rdAddr_1 ? lvtReg_756 : _GEN_5875; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5877 = 10'h2f5 == io_rdAddr_1 ? lvtReg_757 : _GEN_5876; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5878 = 10'h2f6 == io_rdAddr_1 ? lvtReg_758 : _GEN_5877; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5879 = 10'h2f7 == io_rdAddr_1 ? lvtReg_759 : _GEN_5878; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5880 = 10'h2f8 == io_rdAddr_1 ? lvtReg_760 : _GEN_5879; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5881 = 10'h2f9 == io_rdAddr_1 ? lvtReg_761 : _GEN_5880; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5882 = 10'h2fa == io_rdAddr_1 ? lvtReg_762 : _GEN_5881; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5883 = 10'h2fb == io_rdAddr_1 ? lvtReg_763 : _GEN_5882; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5884 = 10'h2fc == io_rdAddr_1 ? lvtReg_764 : _GEN_5883; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5885 = 10'h2fd == io_rdAddr_1 ? lvtReg_765 : _GEN_5884; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5886 = 10'h2fe == io_rdAddr_1 ? lvtReg_766 : _GEN_5885; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5887 = 10'h2ff == io_rdAddr_1 ? lvtReg_767 : _GEN_5886; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5888 = 10'h300 == io_rdAddr_1 ? lvtReg_768 : _GEN_5887; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5889 = 10'h301 == io_rdAddr_1 ? lvtReg_769 : _GEN_5888; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5890 = 10'h302 == io_rdAddr_1 ? lvtReg_770 : _GEN_5889; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5891 = 10'h303 == io_rdAddr_1 ? lvtReg_771 : _GEN_5890; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5892 = 10'h304 == io_rdAddr_1 ? lvtReg_772 : _GEN_5891; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5893 = 10'h305 == io_rdAddr_1 ? lvtReg_773 : _GEN_5892; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5894 = 10'h306 == io_rdAddr_1 ? lvtReg_774 : _GEN_5893; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5895 = 10'h307 == io_rdAddr_1 ? lvtReg_775 : _GEN_5894; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5896 = 10'h308 == io_rdAddr_1 ? lvtReg_776 : _GEN_5895; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5897 = 10'h309 == io_rdAddr_1 ? lvtReg_777 : _GEN_5896; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5898 = 10'h30a == io_rdAddr_1 ? lvtReg_778 : _GEN_5897; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5899 = 10'h30b == io_rdAddr_1 ? lvtReg_779 : _GEN_5898; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5900 = 10'h30c == io_rdAddr_1 ? lvtReg_780 : _GEN_5899; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5901 = 10'h30d == io_rdAddr_1 ? lvtReg_781 : _GEN_5900; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5902 = 10'h30e == io_rdAddr_1 ? lvtReg_782 : _GEN_5901; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5903 = 10'h30f == io_rdAddr_1 ? lvtReg_783 : _GEN_5902; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5904 = 10'h310 == io_rdAddr_1 ? lvtReg_784 : _GEN_5903; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5905 = 10'h311 == io_rdAddr_1 ? lvtReg_785 : _GEN_5904; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5906 = 10'h312 == io_rdAddr_1 ? lvtReg_786 : _GEN_5905; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5907 = 10'h313 == io_rdAddr_1 ? lvtReg_787 : _GEN_5906; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5908 = 10'h314 == io_rdAddr_1 ? lvtReg_788 : _GEN_5907; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5909 = 10'h315 == io_rdAddr_1 ? lvtReg_789 : _GEN_5908; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5910 = 10'h316 == io_rdAddr_1 ? lvtReg_790 : _GEN_5909; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5911 = 10'h317 == io_rdAddr_1 ? lvtReg_791 : _GEN_5910; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5912 = 10'h318 == io_rdAddr_1 ? lvtReg_792 : _GEN_5911; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5913 = 10'h319 == io_rdAddr_1 ? lvtReg_793 : _GEN_5912; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5914 = 10'h31a == io_rdAddr_1 ? lvtReg_794 : _GEN_5913; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5915 = 10'h31b == io_rdAddr_1 ? lvtReg_795 : _GEN_5914; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5916 = 10'h31c == io_rdAddr_1 ? lvtReg_796 : _GEN_5915; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5917 = 10'h31d == io_rdAddr_1 ? lvtReg_797 : _GEN_5916; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5918 = 10'h31e == io_rdAddr_1 ? lvtReg_798 : _GEN_5917; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5919 = 10'h31f == io_rdAddr_1 ? lvtReg_799 : _GEN_5918; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5920 = 10'h320 == io_rdAddr_1 ? lvtReg_800 : _GEN_5919; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5921 = 10'h321 == io_rdAddr_1 ? lvtReg_801 : _GEN_5920; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5922 = 10'h322 == io_rdAddr_1 ? lvtReg_802 : _GEN_5921; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5923 = 10'h323 == io_rdAddr_1 ? lvtReg_803 : _GEN_5922; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5924 = 10'h324 == io_rdAddr_1 ? lvtReg_804 : _GEN_5923; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5925 = 10'h325 == io_rdAddr_1 ? lvtReg_805 : _GEN_5924; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5926 = 10'h326 == io_rdAddr_1 ? lvtReg_806 : _GEN_5925; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5927 = 10'h327 == io_rdAddr_1 ? lvtReg_807 : _GEN_5926; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5928 = 10'h328 == io_rdAddr_1 ? lvtReg_808 : _GEN_5927; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5929 = 10'h329 == io_rdAddr_1 ? lvtReg_809 : _GEN_5928; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5930 = 10'h32a == io_rdAddr_1 ? lvtReg_810 : _GEN_5929; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5931 = 10'h32b == io_rdAddr_1 ? lvtReg_811 : _GEN_5930; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5932 = 10'h32c == io_rdAddr_1 ? lvtReg_812 : _GEN_5931; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5933 = 10'h32d == io_rdAddr_1 ? lvtReg_813 : _GEN_5932; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5934 = 10'h32e == io_rdAddr_1 ? lvtReg_814 : _GEN_5933; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5935 = 10'h32f == io_rdAddr_1 ? lvtReg_815 : _GEN_5934; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5936 = 10'h330 == io_rdAddr_1 ? lvtReg_816 : _GEN_5935; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5937 = 10'h331 == io_rdAddr_1 ? lvtReg_817 : _GEN_5936; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5938 = 10'h332 == io_rdAddr_1 ? lvtReg_818 : _GEN_5937; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5939 = 10'h333 == io_rdAddr_1 ? lvtReg_819 : _GEN_5938; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5940 = 10'h334 == io_rdAddr_1 ? lvtReg_820 : _GEN_5939; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5941 = 10'h335 == io_rdAddr_1 ? lvtReg_821 : _GEN_5940; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5942 = 10'h336 == io_rdAddr_1 ? lvtReg_822 : _GEN_5941; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5943 = 10'h337 == io_rdAddr_1 ? lvtReg_823 : _GEN_5942; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5944 = 10'h338 == io_rdAddr_1 ? lvtReg_824 : _GEN_5943; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5945 = 10'h339 == io_rdAddr_1 ? lvtReg_825 : _GEN_5944; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5946 = 10'h33a == io_rdAddr_1 ? lvtReg_826 : _GEN_5945; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5947 = 10'h33b == io_rdAddr_1 ? lvtReg_827 : _GEN_5946; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5948 = 10'h33c == io_rdAddr_1 ? lvtReg_828 : _GEN_5947; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5949 = 10'h33d == io_rdAddr_1 ? lvtReg_829 : _GEN_5948; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5950 = 10'h33e == io_rdAddr_1 ? lvtReg_830 : _GEN_5949; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5951 = 10'h33f == io_rdAddr_1 ? lvtReg_831 : _GEN_5950; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5952 = 10'h340 == io_rdAddr_1 ? lvtReg_832 : _GEN_5951; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5953 = 10'h341 == io_rdAddr_1 ? lvtReg_833 : _GEN_5952; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5954 = 10'h342 == io_rdAddr_1 ? lvtReg_834 : _GEN_5953; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5955 = 10'h343 == io_rdAddr_1 ? lvtReg_835 : _GEN_5954; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5956 = 10'h344 == io_rdAddr_1 ? lvtReg_836 : _GEN_5955; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5957 = 10'h345 == io_rdAddr_1 ? lvtReg_837 : _GEN_5956; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5958 = 10'h346 == io_rdAddr_1 ? lvtReg_838 : _GEN_5957; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5959 = 10'h347 == io_rdAddr_1 ? lvtReg_839 : _GEN_5958; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5960 = 10'h348 == io_rdAddr_1 ? lvtReg_840 : _GEN_5959; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5961 = 10'h349 == io_rdAddr_1 ? lvtReg_841 : _GEN_5960; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5962 = 10'h34a == io_rdAddr_1 ? lvtReg_842 : _GEN_5961; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5963 = 10'h34b == io_rdAddr_1 ? lvtReg_843 : _GEN_5962; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5964 = 10'h34c == io_rdAddr_1 ? lvtReg_844 : _GEN_5963; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5965 = 10'h34d == io_rdAddr_1 ? lvtReg_845 : _GEN_5964; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5966 = 10'h34e == io_rdAddr_1 ? lvtReg_846 : _GEN_5965; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5967 = 10'h34f == io_rdAddr_1 ? lvtReg_847 : _GEN_5966; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5968 = 10'h350 == io_rdAddr_1 ? lvtReg_848 : _GEN_5967; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5969 = 10'h351 == io_rdAddr_1 ? lvtReg_849 : _GEN_5968; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5970 = 10'h352 == io_rdAddr_1 ? lvtReg_850 : _GEN_5969; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5971 = 10'h353 == io_rdAddr_1 ? lvtReg_851 : _GEN_5970; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5972 = 10'h354 == io_rdAddr_1 ? lvtReg_852 : _GEN_5971; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5973 = 10'h355 == io_rdAddr_1 ? lvtReg_853 : _GEN_5972; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5974 = 10'h356 == io_rdAddr_1 ? lvtReg_854 : _GEN_5973; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5975 = 10'h357 == io_rdAddr_1 ? lvtReg_855 : _GEN_5974; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5976 = 10'h358 == io_rdAddr_1 ? lvtReg_856 : _GEN_5975; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5977 = 10'h359 == io_rdAddr_1 ? lvtReg_857 : _GEN_5976; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5978 = 10'h35a == io_rdAddr_1 ? lvtReg_858 : _GEN_5977; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5979 = 10'h35b == io_rdAddr_1 ? lvtReg_859 : _GEN_5978; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5980 = 10'h35c == io_rdAddr_1 ? lvtReg_860 : _GEN_5979; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5981 = 10'h35d == io_rdAddr_1 ? lvtReg_861 : _GEN_5980; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5982 = 10'h35e == io_rdAddr_1 ? lvtReg_862 : _GEN_5981; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5983 = 10'h35f == io_rdAddr_1 ? lvtReg_863 : _GEN_5982; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5984 = 10'h360 == io_rdAddr_1 ? lvtReg_864 : _GEN_5983; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5985 = 10'h361 == io_rdAddr_1 ? lvtReg_865 : _GEN_5984; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5986 = 10'h362 == io_rdAddr_1 ? lvtReg_866 : _GEN_5985; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5987 = 10'h363 == io_rdAddr_1 ? lvtReg_867 : _GEN_5986; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5988 = 10'h364 == io_rdAddr_1 ? lvtReg_868 : _GEN_5987; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5989 = 10'h365 == io_rdAddr_1 ? lvtReg_869 : _GEN_5988; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5990 = 10'h366 == io_rdAddr_1 ? lvtReg_870 : _GEN_5989; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5991 = 10'h367 == io_rdAddr_1 ? lvtReg_871 : _GEN_5990; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5992 = 10'h368 == io_rdAddr_1 ? lvtReg_872 : _GEN_5991; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5993 = 10'h369 == io_rdAddr_1 ? lvtReg_873 : _GEN_5992; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5994 = 10'h36a == io_rdAddr_1 ? lvtReg_874 : _GEN_5993; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5995 = 10'h36b == io_rdAddr_1 ? lvtReg_875 : _GEN_5994; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5996 = 10'h36c == io_rdAddr_1 ? lvtReg_876 : _GEN_5995; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5997 = 10'h36d == io_rdAddr_1 ? lvtReg_877 : _GEN_5996; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5998 = 10'h36e == io_rdAddr_1 ? lvtReg_878 : _GEN_5997; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_5999 = 10'h36f == io_rdAddr_1 ? lvtReg_879 : _GEN_5998; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6000 = 10'h370 == io_rdAddr_1 ? lvtReg_880 : _GEN_5999; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6001 = 10'h371 == io_rdAddr_1 ? lvtReg_881 : _GEN_6000; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6002 = 10'h372 == io_rdAddr_1 ? lvtReg_882 : _GEN_6001; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6003 = 10'h373 == io_rdAddr_1 ? lvtReg_883 : _GEN_6002; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6004 = 10'h374 == io_rdAddr_1 ? lvtReg_884 : _GEN_6003; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6005 = 10'h375 == io_rdAddr_1 ? lvtReg_885 : _GEN_6004; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6006 = 10'h376 == io_rdAddr_1 ? lvtReg_886 : _GEN_6005; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6007 = 10'h377 == io_rdAddr_1 ? lvtReg_887 : _GEN_6006; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6008 = 10'h378 == io_rdAddr_1 ? lvtReg_888 : _GEN_6007; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6009 = 10'h379 == io_rdAddr_1 ? lvtReg_889 : _GEN_6008; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6010 = 10'h37a == io_rdAddr_1 ? lvtReg_890 : _GEN_6009; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6011 = 10'h37b == io_rdAddr_1 ? lvtReg_891 : _GEN_6010; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6012 = 10'h37c == io_rdAddr_1 ? lvtReg_892 : _GEN_6011; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6013 = 10'h37d == io_rdAddr_1 ? lvtReg_893 : _GEN_6012; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6014 = 10'h37e == io_rdAddr_1 ? lvtReg_894 : _GEN_6013; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6015 = 10'h37f == io_rdAddr_1 ? lvtReg_895 : _GEN_6014; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6016 = 10'h380 == io_rdAddr_1 ? lvtReg_896 : _GEN_6015; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6017 = 10'h381 == io_rdAddr_1 ? lvtReg_897 : _GEN_6016; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6018 = 10'h382 == io_rdAddr_1 ? lvtReg_898 : _GEN_6017; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6019 = 10'h383 == io_rdAddr_1 ? lvtReg_899 : _GEN_6018; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6020 = 10'h384 == io_rdAddr_1 ? lvtReg_900 : _GEN_6019; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6021 = 10'h385 == io_rdAddr_1 ? lvtReg_901 : _GEN_6020; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6022 = 10'h386 == io_rdAddr_1 ? lvtReg_902 : _GEN_6021; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6023 = 10'h387 == io_rdAddr_1 ? lvtReg_903 : _GEN_6022; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6024 = 10'h388 == io_rdAddr_1 ? lvtReg_904 : _GEN_6023; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6025 = 10'h389 == io_rdAddr_1 ? lvtReg_905 : _GEN_6024; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6026 = 10'h38a == io_rdAddr_1 ? lvtReg_906 : _GEN_6025; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6027 = 10'h38b == io_rdAddr_1 ? lvtReg_907 : _GEN_6026; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6028 = 10'h38c == io_rdAddr_1 ? lvtReg_908 : _GEN_6027; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6029 = 10'h38d == io_rdAddr_1 ? lvtReg_909 : _GEN_6028; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6030 = 10'h38e == io_rdAddr_1 ? lvtReg_910 : _GEN_6029; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6031 = 10'h38f == io_rdAddr_1 ? lvtReg_911 : _GEN_6030; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6032 = 10'h390 == io_rdAddr_1 ? lvtReg_912 : _GEN_6031; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6033 = 10'h391 == io_rdAddr_1 ? lvtReg_913 : _GEN_6032; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6034 = 10'h392 == io_rdAddr_1 ? lvtReg_914 : _GEN_6033; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6035 = 10'h393 == io_rdAddr_1 ? lvtReg_915 : _GEN_6034; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6036 = 10'h394 == io_rdAddr_1 ? lvtReg_916 : _GEN_6035; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6037 = 10'h395 == io_rdAddr_1 ? lvtReg_917 : _GEN_6036; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6038 = 10'h396 == io_rdAddr_1 ? lvtReg_918 : _GEN_6037; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6039 = 10'h397 == io_rdAddr_1 ? lvtReg_919 : _GEN_6038; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6040 = 10'h398 == io_rdAddr_1 ? lvtReg_920 : _GEN_6039; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6041 = 10'h399 == io_rdAddr_1 ? lvtReg_921 : _GEN_6040; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6042 = 10'h39a == io_rdAddr_1 ? lvtReg_922 : _GEN_6041; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6043 = 10'h39b == io_rdAddr_1 ? lvtReg_923 : _GEN_6042; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6044 = 10'h39c == io_rdAddr_1 ? lvtReg_924 : _GEN_6043; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6045 = 10'h39d == io_rdAddr_1 ? lvtReg_925 : _GEN_6044; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6046 = 10'h39e == io_rdAddr_1 ? lvtReg_926 : _GEN_6045; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6047 = 10'h39f == io_rdAddr_1 ? lvtReg_927 : _GEN_6046; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6048 = 10'h3a0 == io_rdAddr_1 ? lvtReg_928 : _GEN_6047; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6049 = 10'h3a1 == io_rdAddr_1 ? lvtReg_929 : _GEN_6048; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6050 = 10'h3a2 == io_rdAddr_1 ? lvtReg_930 : _GEN_6049; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6051 = 10'h3a3 == io_rdAddr_1 ? lvtReg_931 : _GEN_6050; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6052 = 10'h3a4 == io_rdAddr_1 ? lvtReg_932 : _GEN_6051; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6053 = 10'h3a5 == io_rdAddr_1 ? lvtReg_933 : _GEN_6052; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6054 = 10'h3a6 == io_rdAddr_1 ? lvtReg_934 : _GEN_6053; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6055 = 10'h3a7 == io_rdAddr_1 ? lvtReg_935 : _GEN_6054; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6056 = 10'h3a8 == io_rdAddr_1 ? lvtReg_936 : _GEN_6055; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6057 = 10'h3a9 == io_rdAddr_1 ? lvtReg_937 : _GEN_6056; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6058 = 10'h3aa == io_rdAddr_1 ? lvtReg_938 : _GEN_6057; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6059 = 10'h3ab == io_rdAddr_1 ? lvtReg_939 : _GEN_6058; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6060 = 10'h3ac == io_rdAddr_1 ? lvtReg_940 : _GEN_6059; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6061 = 10'h3ad == io_rdAddr_1 ? lvtReg_941 : _GEN_6060; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6062 = 10'h3ae == io_rdAddr_1 ? lvtReg_942 : _GEN_6061; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6063 = 10'h3af == io_rdAddr_1 ? lvtReg_943 : _GEN_6062; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6064 = 10'h3b0 == io_rdAddr_1 ? lvtReg_944 : _GEN_6063; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6065 = 10'h3b1 == io_rdAddr_1 ? lvtReg_945 : _GEN_6064; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6066 = 10'h3b2 == io_rdAddr_1 ? lvtReg_946 : _GEN_6065; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6067 = 10'h3b3 == io_rdAddr_1 ? lvtReg_947 : _GEN_6066; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6068 = 10'h3b4 == io_rdAddr_1 ? lvtReg_948 : _GEN_6067; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6069 = 10'h3b5 == io_rdAddr_1 ? lvtReg_949 : _GEN_6068; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6070 = 10'h3b6 == io_rdAddr_1 ? lvtReg_950 : _GEN_6069; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6071 = 10'h3b7 == io_rdAddr_1 ? lvtReg_951 : _GEN_6070; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6072 = 10'h3b8 == io_rdAddr_1 ? lvtReg_952 : _GEN_6071; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6073 = 10'h3b9 == io_rdAddr_1 ? lvtReg_953 : _GEN_6072; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6074 = 10'h3ba == io_rdAddr_1 ? lvtReg_954 : _GEN_6073; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6075 = 10'h3bb == io_rdAddr_1 ? lvtReg_955 : _GEN_6074; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6076 = 10'h3bc == io_rdAddr_1 ? lvtReg_956 : _GEN_6075; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6077 = 10'h3bd == io_rdAddr_1 ? lvtReg_957 : _GEN_6076; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6078 = 10'h3be == io_rdAddr_1 ? lvtReg_958 : _GEN_6077; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6079 = 10'h3bf == io_rdAddr_1 ? lvtReg_959 : _GEN_6078; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6080 = 10'h3c0 == io_rdAddr_1 ? lvtReg_960 : _GEN_6079; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6081 = 10'h3c1 == io_rdAddr_1 ? lvtReg_961 : _GEN_6080; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6082 = 10'h3c2 == io_rdAddr_1 ? lvtReg_962 : _GEN_6081; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6083 = 10'h3c3 == io_rdAddr_1 ? lvtReg_963 : _GEN_6082; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6084 = 10'h3c4 == io_rdAddr_1 ? lvtReg_964 : _GEN_6083; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6085 = 10'h3c5 == io_rdAddr_1 ? lvtReg_965 : _GEN_6084; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6086 = 10'h3c6 == io_rdAddr_1 ? lvtReg_966 : _GEN_6085; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6087 = 10'h3c7 == io_rdAddr_1 ? lvtReg_967 : _GEN_6086; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6088 = 10'h3c8 == io_rdAddr_1 ? lvtReg_968 : _GEN_6087; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6089 = 10'h3c9 == io_rdAddr_1 ? lvtReg_969 : _GEN_6088; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6090 = 10'h3ca == io_rdAddr_1 ? lvtReg_970 : _GEN_6089; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6091 = 10'h3cb == io_rdAddr_1 ? lvtReg_971 : _GEN_6090; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6092 = 10'h3cc == io_rdAddr_1 ? lvtReg_972 : _GEN_6091; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6093 = 10'h3cd == io_rdAddr_1 ? lvtReg_973 : _GEN_6092; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6094 = 10'h3ce == io_rdAddr_1 ? lvtReg_974 : _GEN_6093; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6095 = 10'h3cf == io_rdAddr_1 ? lvtReg_975 : _GEN_6094; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6096 = 10'h3d0 == io_rdAddr_1 ? lvtReg_976 : _GEN_6095; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6097 = 10'h3d1 == io_rdAddr_1 ? lvtReg_977 : _GEN_6096; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6098 = 10'h3d2 == io_rdAddr_1 ? lvtReg_978 : _GEN_6097; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6099 = 10'h3d3 == io_rdAddr_1 ? lvtReg_979 : _GEN_6098; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6100 = 10'h3d4 == io_rdAddr_1 ? lvtReg_980 : _GEN_6099; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6101 = 10'h3d5 == io_rdAddr_1 ? lvtReg_981 : _GEN_6100; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6102 = 10'h3d6 == io_rdAddr_1 ? lvtReg_982 : _GEN_6101; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6103 = 10'h3d7 == io_rdAddr_1 ? lvtReg_983 : _GEN_6102; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6104 = 10'h3d8 == io_rdAddr_1 ? lvtReg_984 : _GEN_6103; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6105 = 10'h3d9 == io_rdAddr_1 ? lvtReg_985 : _GEN_6104; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6106 = 10'h3da == io_rdAddr_1 ? lvtReg_986 : _GEN_6105; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6107 = 10'h3db == io_rdAddr_1 ? lvtReg_987 : _GEN_6106; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6108 = 10'h3dc == io_rdAddr_1 ? lvtReg_988 : _GEN_6107; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6109 = 10'h3dd == io_rdAddr_1 ? lvtReg_989 : _GEN_6108; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6110 = 10'h3de == io_rdAddr_1 ? lvtReg_990 : _GEN_6109; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6111 = 10'h3df == io_rdAddr_1 ? lvtReg_991 : _GEN_6110; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6112 = 10'h3e0 == io_rdAddr_1 ? lvtReg_992 : _GEN_6111; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6113 = 10'h3e1 == io_rdAddr_1 ? lvtReg_993 : _GEN_6112; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6114 = 10'h3e2 == io_rdAddr_1 ? lvtReg_994 : _GEN_6113; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6115 = 10'h3e3 == io_rdAddr_1 ? lvtReg_995 : _GEN_6114; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6116 = 10'h3e4 == io_rdAddr_1 ? lvtReg_996 : _GEN_6115; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6117 = 10'h3e5 == io_rdAddr_1 ? lvtReg_997 : _GEN_6116; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6118 = 10'h3e6 == io_rdAddr_1 ? lvtReg_998 : _GEN_6117; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6119 = 10'h3e7 == io_rdAddr_1 ? lvtReg_999 : _GEN_6118; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6120 = 10'h3e8 == io_rdAddr_1 ? lvtReg_1000 : _GEN_6119; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6121 = 10'h3e9 == io_rdAddr_1 ? lvtReg_1001 : _GEN_6120; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6122 = 10'h3ea == io_rdAddr_1 ? lvtReg_1002 : _GEN_6121; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6123 = 10'h3eb == io_rdAddr_1 ? lvtReg_1003 : _GEN_6122; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6124 = 10'h3ec == io_rdAddr_1 ? lvtReg_1004 : _GEN_6123; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6125 = 10'h3ed == io_rdAddr_1 ? lvtReg_1005 : _GEN_6124; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6126 = 10'h3ee == io_rdAddr_1 ? lvtReg_1006 : _GEN_6125; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6127 = 10'h3ef == io_rdAddr_1 ? lvtReg_1007 : _GEN_6126; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6128 = 10'h3f0 == io_rdAddr_1 ? lvtReg_1008 : _GEN_6127; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6129 = 10'h3f1 == io_rdAddr_1 ? lvtReg_1009 : _GEN_6128; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6130 = 10'h3f2 == io_rdAddr_1 ? lvtReg_1010 : _GEN_6129; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6131 = 10'h3f3 == io_rdAddr_1 ? lvtReg_1011 : _GEN_6130; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6132 = 10'h3f4 == io_rdAddr_1 ? lvtReg_1012 : _GEN_6131; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6133 = 10'h3f5 == io_rdAddr_1 ? lvtReg_1013 : _GEN_6132; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6134 = 10'h3f6 == io_rdAddr_1 ? lvtReg_1014 : _GEN_6133; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6135 = 10'h3f7 == io_rdAddr_1 ? lvtReg_1015 : _GEN_6134; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6136 = 10'h3f8 == io_rdAddr_1 ? lvtReg_1016 : _GEN_6135; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6137 = 10'h3f9 == io_rdAddr_1 ? lvtReg_1017 : _GEN_6136; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6138 = 10'h3fa == io_rdAddr_1 ? lvtReg_1018 : _GEN_6137; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6139 = 10'h3fb == io_rdAddr_1 ? lvtReg_1019 : _GEN_6138; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6140 = 10'h3fc == io_rdAddr_1 ? lvtReg_1020 : _GEN_6139; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6141 = 10'h3fd == io_rdAddr_1 ? lvtReg_1021 : _GEN_6140; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_6142 = 10'h3fe == io_rdAddr_1 ? lvtReg_1022 : _GEN_6141; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_0 = 10'h3ff == io_rdAddr_0 ? lvtReg_1023 : _GEN_5118; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_1 = 10'h3ff == io_rdAddr_1 ? lvtReg_1023 : _GEN_6142; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  always @(posedge clock) begin
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_0 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_0 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_0 <= _GEN_1024;
      end
    end else begin
      lvtReg_0 <= _GEN_1024;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1 <= _GEN_1025;
      end
    end else begin
      lvtReg_1 <= _GEN_1025;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_2 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_2 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_2 <= _GEN_1026;
      end
    end else begin
      lvtReg_2 <= _GEN_1026;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_3 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_3 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_3 <= _GEN_1027;
      end
    end else begin
      lvtReg_3 <= _GEN_1027;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_4 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_4 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_4 <= _GEN_1028;
      end
    end else begin
      lvtReg_4 <= _GEN_1028;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_5 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_5 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_5 <= _GEN_1029;
      end
    end else begin
      lvtReg_5 <= _GEN_1029;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_6 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_6 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_6 <= _GEN_1030;
      end
    end else begin
      lvtReg_6 <= _GEN_1030;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_7 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_7 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_7 <= _GEN_1031;
      end
    end else begin
      lvtReg_7 <= _GEN_1031;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_8 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_8 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_8 <= _GEN_1032;
      end
    end else begin
      lvtReg_8 <= _GEN_1032;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_9 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_9 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_9 <= _GEN_1033;
      end
    end else begin
      lvtReg_9 <= _GEN_1033;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_10 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_10 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_10 <= _GEN_1034;
      end
    end else begin
      lvtReg_10 <= _GEN_1034;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_11 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_11 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_11 <= _GEN_1035;
      end
    end else begin
      lvtReg_11 <= _GEN_1035;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_12 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_12 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_12 <= _GEN_1036;
      end
    end else begin
      lvtReg_12 <= _GEN_1036;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_13 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_13 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_13 <= _GEN_1037;
      end
    end else begin
      lvtReg_13 <= _GEN_1037;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_14 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_14 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_14 <= _GEN_1038;
      end
    end else begin
      lvtReg_14 <= _GEN_1038;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_15 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_15 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_15 <= _GEN_1039;
      end
    end else begin
      lvtReg_15 <= _GEN_1039;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_16 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_16 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_16 <= _GEN_1040;
      end
    end else begin
      lvtReg_16 <= _GEN_1040;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_17 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_17 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_17 <= _GEN_1041;
      end
    end else begin
      lvtReg_17 <= _GEN_1041;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_18 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_18 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_18 <= _GEN_1042;
      end
    end else begin
      lvtReg_18 <= _GEN_1042;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_19 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_19 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_19 <= _GEN_1043;
      end
    end else begin
      lvtReg_19 <= _GEN_1043;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_20 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_20 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_20 <= _GEN_1044;
      end
    end else begin
      lvtReg_20 <= _GEN_1044;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_21 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_21 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_21 <= _GEN_1045;
      end
    end else begin
      lvtReg_21 <= _GEN_1045;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_22 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_22 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_22 <= _GEN_1046;
      end
    end else begin
      lvtReg_22 <= _GEN_1046;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_23 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_23 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_23 <= _GEN_1047;
      end
    end else begin
      lvtReg_23 <= _GEN_1047;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_24 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_24 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_24 <= _GEN_1048;
      end
    end else begin
      lvtReg_24 <= _GEN_1048;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_25 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_25 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_25 <= _GEN_1049;
      end
    end else begin
      lvtReg_25 <= _GEN_1049;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_26 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_26 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_26 <= _GEN_1050;
      end
    end else begin
      lvtReg_26 <= _GEN_1050;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_27 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_27 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_27 <= _GEN_1051;
      end
    end else begin
      lvtReg_27 <= _GEN_1051;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_28 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_28 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_28 <= _GEN_1052;
      end
    end else begin
      lvtReg_28 <= _GEN_1052;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_29 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_29 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_29 <= _GEN_1053;
      end
    end else begin
      lvtReg_29 <= _GEN_1053;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_30 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_30 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_30 <= _GEN_1054;
      end
    end else begin
      lvtReg_30 <= _GEN_1054;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_31 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_31 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_31 <= _GEN_1055;
      end
    end else begin
      lvtReg_31 <= _GEN_1055;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_32 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_32 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_32 <= _GEN_1056;
      end
    end else begin
      lvtReg_32 <= _GEN_1056;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_33 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_33 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_33 <= _GEN_1057;
      end
    end else begin
      lvtReg_33 <= _GEN_1057;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_34 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_34 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_34 <= _GEN_1058;
      end
    end else begin
      lvtReg_34 <= _GEN_1058;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_35 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_35 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_35 <= _GEN_1059;
      end
    end else begin
      lvtReg_35 <= _GEN_1059;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_36 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_36 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_36 <= _GEN_1060;
      end
    end else begin
      lvtReg_36 <= _GEN_1060;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_37 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_37 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_37 <= _GEN_1061;
      end
    end else begin
      lvtReg_37 <= _GEN_1061;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_38 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_38 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_38 <= _GEN_1062;
      end
    end else begin
      lvtReg_38 <= _GEN_1062;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_39 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_39 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_39 <= _GEN_1063;
      end
    end else begin
      lvtReg_39 <= _GEN_1063;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_40 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_40 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_40 <= _GEN_1064;
      end
    end else begin
      lvtReg_40 <= _GEN_1064;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_41 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_41 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_41 <= _GEN_1065;
      end
    end else begin
      lvtReg_41 <= _GEN_1065;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_42 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_42 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_42 <= _GEN_1066;
      end
    end else begin
      lvtReg_42 <= _GEN_1066;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_43 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_43 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_43 <= _GEN_1067;
      end
    end else begin
      lvtReg_43 <= _GEN_1067;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_44 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_44 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_44 <= _GEN_1068;
      end
    end else begin
      lvtReg_44 <= _GEN_1068;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_45 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_45 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_45 <= _GEN_1069;
      end
    end else begin
      lvtReg_45 <= _GEN_1069;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_46 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_46 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_46 <= _GEN_1070;
      end
    end else begin
      lvtReg_46 <= _GEN_1070;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_47 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_47 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_47 <= _GEN_1071;
      end
    end else begin
      lvtReg_47 <= _GEN_1071;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_48 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_48 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_48 <= _GEN_1072;
      end
    end else begin
      lvtReg_48 <= _GEN_1072;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_49 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_49 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_49 <= _GEN_1073;
      end
    end else begin
      lvtReg_49 <= _GEN_1073;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_50 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_50 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_50 <= _GEN_1074;
      end
    end else begin
      lvtReg_50 <= _GEN_1074;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_51 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_51 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_51 <= _GEN_1075;
      end
    end else begin
      lvtReg_51 <= _GEN_1075;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_52 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_52 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_52 <= _GEN_1076;
      end
    end else begin
      lvtReg_52 <= _GEN_1076;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_53 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_53 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_53 <= _GEN_1077;
      end
    end else begin
      lvtReg_53 <= _GEN_1077;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_54 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_54 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_54 <= _GEN_1078;
      end
    end else begin
      lvtReg_54 <= _GEN_1078;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_55 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_55 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_55 <= _GEN_1079;
      end
    end else begin
      lvtReg_55 <= _GEN_1079;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_56 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_56 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_56 <= _GEN_1080;
      end
    end else begin
      lvtReg_56 <= _GEN_1080;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_57 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_57 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_57 <= _GEN_1081;
      end
    end else begin
      lvtReg_57 <= _GEN_1081;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_58 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_58 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_58 <= _GEN_1082;
      end
    end else begin
      lvtReg_58 <= _GEN_1082;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_59 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_59 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_59 <= _GEN_1083;
      end
    end else begin
      lvtReg_59 <= _GEN_1083;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_60 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_60 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_60 <= _GEN_1084;
      end
    end else begin
      lvtReg_60 <= _GEN_1084;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_61 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_61 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_61 <= _GEN_1085;
      end
    end else begin
      lvtReg_61 <= _GEN_1085;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_62 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_62 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_62 <= _GEN_1086;
      end
    end else begin
      lvtReg_62 <= _GEN_1086;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_63 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_63 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_63 <= _GEN_1087;
      end
    end else begin
      lvtReg_63 <= _GEN_1087;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_64 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h40 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_64 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_64 <= _GEN_1088;
      end
    end else begin
      lvtReg_64 <= _GEN_1088;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_65 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h41 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_65 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_65 <= _GEN_1089;
      end
    end else begin
      lvtReg_65 <= _GEN_1089;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_66 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h42 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_66 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_66 <= _GEN_1090;
      end
    end else begin
      lvtReg_66 <= _GEN_1090;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_67 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h43 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_67 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_67 <= _GEN_1091;
      end
    end else begin
      lvtReg_67 <= _GEN_1091;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_68 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h44 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_68 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_68 <= _GEN_1092;
      end
    end else begin
      lvtReg_68 <= _GEN_1092;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_69 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h45 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_69 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_69 <= _GEN_1093;
      end
    end else begin
      lvtReg_69 <= _GEN_1093;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_70 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h46 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_70 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_70 <= _GEN_1094;
      end
    end else begin
      lvtReg_70 <= _GEN_1094;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_71 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h47 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_71 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_71 <= _GEN_1095;
      end
    end else begin
      lvtReg_71 <= _GEN_1095;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_72 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h48 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_72 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_72 <= _GEN_1096;
      end
    end else begin
      lvtReg_72 <= _GEN_1096;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_73 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h49 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_73 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_73 <= _GEN_1097;
      end
    end else begin
      lvtReg_73 <= _GEN_1097;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_74 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_74 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_74 <= _GEN_1098;
      end
    end else begin
      lvtReg_74 <= _GEN_1098;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_75 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_75 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_75 <= _GEN_1099;
      end
    end else begin
      lvtReg_75 <= _GEN_1099;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_76 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_76 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_76 <= _GEN_1100;
      end
    end else begin
      lvtReg_76 <= _GEN_1100;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_77 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_77 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_77 <= _GEN_1101;
      end
    end else begin
      lvtReg_77 <= _GEN_1101;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_78 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_78 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_78 <= _GEN_1102;
      end
    end else begin
      lvtReg_78 <= _GEN_1102;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_79 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h4f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_79 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_79 <= _GEN_1103;
      end
    end else begin
      lvtReg_79 <= _GEN_1103;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_80 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h50 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_80 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_80 <= _GEN_1104;
      end
    end else begin
      lvtReg_80 <= _GEN_1104;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_81 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h51 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_81 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_81 <= _GEN_1105;
      end
    end else begin
      lvtReg_81 <= _GEN_1105;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_82 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h52 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_82 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_82 <= _GEN_1106;
      end
    end else begin
      lvtReg_82 <= _GEN_1106;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_83 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h53 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_83 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_83 <= _GEN_1107;
      end
    end else begin
      lvtReg_83 <= _GEN_1107;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_84 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h54 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_84 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_84 <= _GEN_1108;
      end
    end else begin
      lvtReg_84 <= _GEN_1108;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_85 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h55 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_85 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_85 <= _GEN_1109;
      end
    end else begin
      lvtReg_85 <= _GEN_1109;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_86 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h56 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_86 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_86 <= _GEN_1110;
      end
    end else begin
      lvtReg_86 <= _GEN_1110;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_87 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h57 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_87 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_87 <= _GEN_1111;
      end
    end else begin
      lvtReg_87 <= _GEN_1111;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_88 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h58 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_88 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_88 <= _GEN_1112;
      end
    end else begin
      lvtReg_88 <= _GEN_1112;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_89 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h59 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_89 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_89 <= _GEN_1113;
      end
    end else begin
      lvtReg_89 <= _GEN_1113;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_90 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_90 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_90 <= _GEN_1114;
      end
    end else begin
      lvtReg_90 <= _GEN_1114;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_91 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_91 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_91 <= _GEN_1115;
      end
    end else begin
      lvtReg_91 <= _GEN_1115;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_92 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_92 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_92 <= _GEN_1116;
      end
    end else begin
      lvtReg_92 <= _GEN_1116;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_93 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_93 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_93 <= _GEN_1117;
      end
    end else begin
      lvtReg_93 <= _GEN_1117;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_94 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_94 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_94 <= _GEN_1118;
      end
    end else begin
      lvtReg_94 <= _GEN_1118;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_95 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h5f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_95 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_95 <= _GEN_1119;
      end
    end else begin
      lvtReg_95 <= _GEN_1119;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_96 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h60 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_96 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_96 <= _GEN_1120;
      end
    end else begin
      lvtReg_96 <= _GEN_1120;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_97 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h61 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_97 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_97 <= _GEN_1121;
      end
    end else begin
      lvtReg_97 <= _GEN_1121;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_98 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h62 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_98 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_98 <= _GEN_1122;
      end
    end else begin
      lvtReg_98 <= _GEN_1122;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_99 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h63 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_99 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_99 <= _GEN_1123;
      end
    end else begin
      lvtReg_99 <= _GEN_1123;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_100 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h64 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_100 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_100 <= _GEN_1124;
      end
    end else begin
      lvtReg_100 <= _GEN_1124;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_101 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h65 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_101 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_101 <= _GEN_1125;
      end
    end else begin
      lvtReg_101 <= _GEN_1125;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_102 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h66 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_102 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_102 <= _GEN_1126;
      end
    end else begin
      lvtReg_102 <= _GEN_1126;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_103 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h67 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_103 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_103 <= _GEN_1127;
      end
    end else begin
      lvtReg_103 <= _GEN_1127;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_104 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h68 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_104 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_104 <= _GEN_1128;
      end
    end else begin
      lvtReg_104 <= _GEN_1128;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_105 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h69 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_105 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_105 <= _GEN_1129;
      end
    end else begin
      lvtReg_105 <= _GEN_1129;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_106 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_106 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_106 <= _GEN_1130;
      end
    end else begin
      lvtReg_106 <= _GEN_1130;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_107 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_107 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_107 <= _GEN_1131;
      end
    end else begin
      lvtReg_107 <= _GEN_1131;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_108 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_108 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_108 <= _GEN_1132;
      end
    end else begin
      lvtReg_108 <= _GEN_1132;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_109 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_109 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_109 <= _GEN_1133;
      end
    end else begin
      lvtReg_109 <= _GEN_1133;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_110 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_110 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_110 <= _GEN_1134;
      end
    end else begin
      lvtReg_110 <= _GEN_1134;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_111 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h6f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_111 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_111 <= _GEN_1135;
      end
    end else begin
      lvtReg_111 <= _GEN_1135;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_112 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h70 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_112 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_112 <= _GEN_1136;
      end
    end else begin
      lvtReg_112 <= _GEN_1136;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_113 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h71 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_113 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_113 <= _GEN_1137;
      end
    end else begin
      lvtReg_113 <= _GEN_1137;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_114 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h72 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_114 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_114 <= _GEN_1138;
      end
    end else begin
      lvtReg_114 <= _GEN_1138;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_115 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h73 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_115 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_115 <= _GEN_1139;
      end
    end else begin
      lvtReg_115 <= _GEN_1139;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_116 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h74 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_116 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_116 <= _GEN_1140;
      end
    end else begin
      lvtReg_116 <= _GEN_1140;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_117 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h75 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_117 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_117 <= _GEN_1141;
      end
    end else begin
      lvtReg_117 <= _GEN_1141;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_118 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h76 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_118 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_118 <= _GEN_1142;
      end
    end else begin
      lvtReg_118 <= _GEN_1142;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_119 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h77 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_119 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_119 <= _GEN_1143;
      end
    end else begin
      lvtReg_119 <= _GEN_1143;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_120 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h78 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_120 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_120 <= _GEN_1144;
      end
    end else begin
      lvtReg_120 <= _GEN_1144;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_121 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h79 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_121 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_121 <= _GEN_1145;
      end
    end else begin
      lvtReg_121 <= _GEN_1145;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_122 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_122 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_122 <= _GEN_1146;
      end
    end else begin
      lvtReg_122 <= _GEN_1146;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_123 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_123 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_123 <= _GEN_1147;
      end
    end else begin
      lvtReg_123 <= _GEN_1147;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_124 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_124 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_124 <= _GEN_1148;
      end
    end else begin
      lvtReg_124 <= _GEN_1148;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_125 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_125 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_125 <= _GEN_1149;
      end
    end else begin
      lvtReg_125 <= _GEN_1149;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_126 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_126 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_126 <= _GEN_1150;
      end
    end else begin
      lvtReg_126 <= _GEN_1150;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_127 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h7f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_127 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_127 <= _GEN_1151;
      end
    end else begin
      lvtReg_127 <= _GEN_1151;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_128 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h80 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_128 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_128 <= _GEN_1152;
      end
    end else begin
      lvtReg_128 <= _GEN_1152;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_129 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h81 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_129 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_129 <= _GEN_1153;
      end
    end else begin
      lvtReg_129 <= _GEN_1153;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_130 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h82 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_130 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_130 <= _GEN_1154;
      end
    end else begin
      lvtReg_130 <= _GEN_1154;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_131 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h83 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_131 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_131 <= _GEN_1155;
      end
    end else begin
      lvtReg_131 <= _GEN_1155;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_132 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h84 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_132 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_132 <= _GEN_1156;
      end
    end else begin
      lvtReg_132 <= _GEN_1156;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_133 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h85 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_133 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_133 <= _GEN_1157;
      end
    end else begin
      lvtReg_133 <= _GEN_1157;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_134 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h86 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_134 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_134 <= _GEN_1158;
      end
    end else begin
      lvtReg_134 <= _GEN_1158;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_135 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h87 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_135 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_135 <= _GEN_1159;
      end
    end else begin
      lvtReg_135 <= _GEN_1159;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_136 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h88 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_136 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_136 <= _GEN_1160;
      end
    end else begin
      lvtReg_136 <= _GEN_1160;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_137 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h89 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_137 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_137 <= _GEN_1161;
      end
    end else begin
      lvtReg_137 <= _GEN_1161;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_138 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_138 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_138 <= _GEN_1162;
      end
    end else begin
      lvtReg_138 <= _GEN_1162;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_139 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_139 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_139 <= _GEN_1163;
      end
    end else begin
      lvtReg_139 <= _GEN_1163;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_140 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_140 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_140 <= _GEN_1164;
      end
    end else begin
      lvtReg_140 <= _GEN_1164;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_141 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_141 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_141 <= _GEN_1165;
      end
    end else begin
      lvtReg_141 <= _GEN_1165;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_142 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_142 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_142 <= _GEN_1166;
      end
    end else begin
      lvtReg_142 <= _GEN_1166;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_143 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h8f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_143 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_143 <= _GEN_1167;
      end
    end else begin
      lvtReg_143 <= _GEN_1167;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_144 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h90 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_144 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_144 <= _GEN_1168;
      end
    end else begin
      lvtReg_144 <= _GEN_1168;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_145 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h91 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_145 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_145 <= _GEN_1169;
      end
    end else begin
      lvtReg_145 <= _GEN_1169;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_146 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h92 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_146 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_146 <= _GEN_1170;
      end
    end else begin
      lvtReg_146 <= _GEN_1170;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_147 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h93 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_147 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_147 <= _GEN_1171;
      end
    end else begin
      lvtReg_147 <= _GEN_1171;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_148 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h94 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_148 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_148 <= _GEN_1172;
      end
    end else begin
      lvtReg_148 <= _GEN_1172;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_149 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h95 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_149 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_149 <= _GEN_1173;
      end
    end else begin
      lvtReg_149 <= _GEN_1173;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_150 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h96 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_150 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_150 <= _GEN_1174;
      end
    end else begin
      lvtReg_150 <= _GEN_1174;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_151 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h97 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_151 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_151 <= _GEN_1175;
      end
    end else begin
      lvtReg_151 <= _GEN_1175;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_152 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h98 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_152 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_152 <= _GEN_1176;
      end
    end else begin
      lvtReg_152 <= _GEN_1176;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_153 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h99 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_153 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_153 <= _GEN_1177;
      end
    end else begin
      lvtReg_153 <= _GEN_1177;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_154 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_154 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_154 <= _GEN_1178;
      end
    end else begin
      lvtReg_154 <= _GEN_1178;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_155 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_155 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_155 <= _GEN_1179;
      end
    end else begin
      lvtReg_155 <= _GEN_1179;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_156 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_156 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_156 <= _GEN_1180;
      end
    end else begin
      lvtReg_156 <= _GEN_1180;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_157 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_157 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_157 <= _GEN_1181;
      end
    end else begin
      lvtReg_157 <= _GEN_1181;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_158 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_158 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_158 <= _GEN_1182;
      end
    end else begin
      lvtReg_158 <= _GEN_1182;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_159 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h9f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_159 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_159 <= _GEN_1183;
      end
    end else begin
      lvtReg_159 <= _GEN_1183;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_160 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_160 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_160 <= _GEN_1184;
      end
    end else begin
      lvtReg_160 <= _GEN_1184;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_161 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_161 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_161 <= _GEN_1185;
      end
    end else begin
      lvtReg_161 <= _GEN_1185;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_162 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_162 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_162 <= _GEN_1186;
      end
    end else begin
      lvtReg_162 <= _GEN_1186;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_163 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_163 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_163 <= _GEN_1187;
      end
    end else begin
      lvtReg_163 <= _GEN_1187;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_164 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_164 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_164 <= _GEN_1188;
      end
    end else begin
      lvtReg_164 <= _GEN_1188;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_165 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_165 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_165 <= _GEN_1189;
      end
    end else begin
      lvtReg_165 <= _GEN_1189;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_166 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_166 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_166 <= _GEN_1190;
      end
    end else begin
      lvtReg_166 <= _GEN_1190;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_167 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_167 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_167 <= _GEN_1191;
      end
    end else begin
      lvtReg_167 <= _GEN_1191;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_168 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_168 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_168 <= _GEN_1192;
      end
    end else begin
      lvtReg_168 <= _GEN_1192;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_169 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'ha9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_169 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_169 <= _GEN_1193;
      end
    end else begin
      lvtReg_169 <= _GEN_1193;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_170 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'haa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_170 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_170 <= _GEN_1194;
      end
    end else begin
      lvtReg_170 <= _GEN_1194;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_171 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hab == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_171 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_171 <= _GEN_1195;
      end
    end else begin
      lvtReg_171 <= _GEN_1195;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_172 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hac == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_172 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_172 <= _GEN_1196;
      end
    end else begin
      lvtReg_172 <= _GEN_1196;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_173 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'had == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_173 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_173 <= _GEN_1197;
      end
    end else begin
      lvtReg_173 <= _GEN_1197;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_174 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hae == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_174 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_174 <= _GEN_1198;
      end
    end else begin
      lvtReg_174 <= _GEN_1198;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_175 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'haf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_175 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_175 <= _GEN_1199;
      end
    end else begin
      lvtReg_175 <= _GEN_1199;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_176 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_176 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_176 <= _GEN_1200;
      end
    end else begin
      lvtReg_176 <= _GEN_1200;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_177 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_177 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_177 <= _GEN_1201;
      end
    end else begin
      lvtReg_177 <= _GEN_1201;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_178 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_178 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_178 <= _GEN_1202;
      end
    end else begin
      lvtReg_178 <= _GEN_1202;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_179 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_179 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_179 <= _GEN_1203;
      end
    end else begin
      lvtReg_179 <= _GEN_1203;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_180 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_180 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_180 <= _GEN_1204;
      end
    end else begin
      lvtReg_180 <= _GEN_1204;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_181 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_181 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_181 <= _GEN_1205;
      end
    end else begin
      lvtReg_181 <= _GEN_1205;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_182 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_182 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_182 <= _GEN_1206;
      end
    end else begin
      lvtReg_182 <= _GEN_1206;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_183 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_183 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_183 <= _GEN_1207;
      end
    end else begin
      lvtReg_183 <= _GEN_1207;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_184 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_184 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_184 <= _GEN_1208;
      end
    end else begin
      lvtReg_184 <= _GEN_1208;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_185 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hb9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_185 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_185 <= _GEN_1209;
      end
    end else begin
      lvtReg_185 <= _GEN_1209;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_186 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hba == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_186 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_186 <= _GEN_1210;
      end
    end else begin
      lvtReg_186 <= _GEN_1210;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_187 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hbb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_187 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_187 <= _GEN_1211;
      end
    end else begin
      lvtReg_187 <= _GEN_1211;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_188 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hbc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_188 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_188 <= _GEN_1212;
      end
    end else begin
      lvtReg_188 <= _GEN_1212;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_189 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hbd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_189 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_189 <= _GEN_1213;
      end
    end else begin
      lvtReg_189 <= _GEN_1213;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_190 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hbe == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_190 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_190 <= _GEN_1214;
      end
    end else begin
      lvtReg_190 <= _GEN_1214;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_191 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hbf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_191 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_191 <= _GEN_1215;
      end
    end else begin
      lvtReg_191 <= _GEN_1215;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_192 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_192 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_192 <= _GEN_1216;
      end
    end else begin
      lvtReg_192 <= _GEN_1216;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_193 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_193 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_193 <= _GEN_1217;
      end
    end else begin
      lvtReg_193 <= _GEN_1217;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_194 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_194 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_194 <= _GEN_1218;
      end
    end else begin
      lvtReg_194 <= _GEN_1218;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_195 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_195 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_195 <= _GEN_1219;
      end
    end else begin
      lvtReg_195 <= _GEN_1219;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_196 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_196 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_196 <= _GEN_1220;
      end
    end else begin
      lvtReg_196 <= _GEN_1220;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_197 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_197 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_197 <= _GEN_1221;
      end
    end else begin
      lvtReg_197 <= _GEN_1221;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_198 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_198 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_198 <= _GEN_1222;
      end
    end else begin
      lvtReg_198 <= _GEN_1222;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_199 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_199 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_199 <= _GEN_1223;
      end
    end else begin
      lvtReg_199 <= _GEN_1223;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_200 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_200 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_200 <= _GEN_1224;
      end
    end else begin
      lvtReg_200 <= _GEN_1224;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_201 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hc9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_201 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_201 <= _GEN_1225;
      end
    end else begin
      lvtReg_201 <= _GEN_1225;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_202 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hca == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_202 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_202 <= _GEN_1226;
      end
    end else begin
      lvtReg_202 <= _GEN_1226;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_203 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hcb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_203 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_203 <= _GEN_1227;
      end
    end else begin
      lvtReg_203 <= _GEN_1227;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_204 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hcc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_204 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_204 <= _GEN_1228;
      end
    end else begin
      lvtReg_204 <= _GEN_1228;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_205 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hcd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_205 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_205 <= _GEN_1229;
      end
    end else begin
      lvtReg_205 <= _GEN_1229;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_206 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hce == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_206 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_206 <= _GEN_1230;
      end
    end else begin
      lvtReg_206 <= _GEN_1230;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_207 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hcf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_207 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_207 <= _GEN_1231;
      end
    end else begin
      lvtReg_207 <= _GEN_1231;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_208 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_208 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_208 <= _GEN_1232;
      end
    end else begin
      lvtReg_208 <= _GEN_1232;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_209 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_209 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_209 <= _GEN_1233;
      end
    end else begin
      lvtReg_209 <= _GEN_1233;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_210 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_210 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_210 <= _GEN_1234;
      end
    end else begin
      lvtReg_210 <= _GEN_1234;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_211 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_211 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_211 <= _GEN_1235;
      end
    end else begin
      lvtReg_211 <= _GEN_1235;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_212 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_212 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_212 <= _GEN_1236;
      end
    end else begin
      lvtReg_212 <= _GEN_1236;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_213 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_213 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_213 <= _GEN_1237;
      end
    end else begin
      lvtReg_213 <= _GEN_1237;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_214 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_214 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_214 <= _GEN_1238;
      end
    end else begin
      lvtReg_214 <= _GEN_1238;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_215 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_215 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_215 <= _GEN_1239;
      end
    end else begin
      lvtReg_215 <= _GEN_1239;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_216 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_216 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_216 <= _GEN_1240;
      end
    end else begin
      lvtReg_216 <= _GEN_1240;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_217 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hd9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_217 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_217 <= _GEN_1241;
      end
    end else begin
      lvtReg_217 <= _GEN_1241;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_218 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hda == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_218 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_218 <= _GEN_1242;
      end
    end else begin
      lvtReg_218 <= _GEN_1242;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_219 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hdb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_219 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_219 <= _GEN_1243;
      end
    end else begin
      lvtReg_219 <= _GEN_1243;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_220 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hdc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_220 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_220 <= _GEN_1244;
      end
    end else begin
      lvtReg_220 <= _GEN_1244;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_221 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hdd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_221 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_221 <= _GEN_1245;
      end
    end else begin
      lvtReg_221 <= _GEN_1245;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_222 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hde == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_222 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_222 <= _GEN_1246;
      end
    end else begin
      lvtReg_222 <= _GEN_1246;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_223 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hdf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_223 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_223 <= _GEN_1247;
      end
    end else begin
      lvtReg_223 <= _GEN_1247;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_224 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_224 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_224 <= _GEN_1248;
      end
    end else begin
      lvtReg_224 <= _GEN_1248;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_225 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_225 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_225 <= _GEN_1249;
      end
    end else begin
      lvtReg_225 <= _GEN_1249;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_226 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_226 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_226 <= _GEN_1250;
      end
    end else begin
      lvtReg_226 <= _GEN_1250;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_227 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_227 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_227 <= _GEN_1251;
      end
    end else begin
      lvtReg_227 <= _GEN_1251;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_228 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_228 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_228 <= _GEN_1252;
      end
    end else begin
      lvtReg_228 <= _GEN_1252;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_229 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_229 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_229 <= _GEN_1253;
      end
    end else begin
      lvtReg_229 <= _GEN_1253;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_230 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_230 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_230 <= _GEN_1254;
      end
    end else begin
      lvtReg_230 <= _GEN_1254;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_231 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_231 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_231 <= _GEN_1255;
      end
    end else begin
      lvtReg_231 <= _GEN_1255;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_232 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_232 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_232 <= _GEN_1256;
      end
    end else begin
      lvtReg_232 <= _GEN_1256;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_233 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'he9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_233 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_233 <= _GEN_1257;
      end
    end else begin
      lvtReg_233 <= _GEN_1257;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_234 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hea == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_234 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_234 <= _GEN_1258;
      end
    end else begin
      lvtReg_234 <= _GEN_1258;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_235 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'heb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_235 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_235 <= _GEN_1259;
      end
    end else begin
      lvtReg_235 <= _GEN_1259;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_236 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hec == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_236 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_236 <= _GEN_1260;
      end
    end else begin
      lvtReg_236 <= _GEN_1260;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_237 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hed == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_237 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_237 <= _GEN_1261;
      end
    end else begin
      lvtReg_237 <= _GEN_1261;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_238 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hee == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_238 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_238 <= _GEN_1262;
      end
    end else begin
      lvtReg_238 <= _GEN_1262;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_239 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hef == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_239 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_239 <= _GEN_1263;
      end
    end else begin
      lvtReg_239 <= _GEN_1263;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_240 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_240 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_240 <= _GEN_1264;
      end
    end else begin
      lvtReg_240 <= _GEN_1264;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_241 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_241 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_241 <= _GEN_1265;
      end
    end else begin
      lvtReg_241 <= _GEN_1265;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_242 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_242 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_242 <= _GEN_1266;
      end
    end else begin
      lvtReg_242 <= _GEN_1266;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_243 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_243 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_243 <= _GEN_1267;
      end
    end else begin
      lvtReg_243 <= _GEN_1267;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_244 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_244 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_244 <= _GEN_1268;
      end
    end else begin
      lvtReg_244 <= _GEN_1268;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_245 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_245 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_245 <= _GEN_1269;
      end
    end else begin
      lvtReg_245 <= _GEN_1269;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_246 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_246 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_246 <= _GEN_1270;
      end
    end else begin
      lvtReg_246 <= _GEN_1270;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_247 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_247 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_247 <= _GEN_1271;
      end
    end else begin
      lvtReg_247 <= _GEN_1271;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_248 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_248 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_248 <= _GEN_1272;
      end
    end else begin
      lvtReg_248 <= _GEN_1272;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_249 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hf9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_249 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_249 <= _GEN_1273;
      end
    end else begin
      lvtReg_249 <= _GEN_1273;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_250 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hfa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_250 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_250 <= _GEN_1274;
      end
    end else begin
      lvtReg_250 <= _GEN_1274;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_251 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hfb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_251 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_251 <= _GEN_1275;
      end
    end else begin
      lvtReg_251 <= _GEN_1275;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_252 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hfc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_252 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_252 <= _GEN_1276;
      end
    end else begin
      lvtReg_252 <= _GEN_1276;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_253 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hfd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_253 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_253 <= _GEN_1277;
      end
    end else begin
      lvtReg_253 <= _GEN_1277;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_254 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hfe == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_254 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_254 <= _GEN_1278;
      end
    end else begin
      lvtReg_254 <= _GEN_1278;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_255 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'hff == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_255 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_255 <= _GEN_1279;
      end
    end else begin
      lvtReg_255 <= _GEN_1279;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_256 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h100 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_256 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_256 <= _GEN_1280;
      end
    end else begin
      lvtReg_256 <= _GEN_1280;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_257 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h101 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_257 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_257 <= _GEN_1281;
      end
    end else begin
      lvtReg_257 <= _GEN_1281;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_258 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h102 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_258 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_258 <= _GEN_1282;
      end
    end else begin
      lvtReg_258 <= _GEN_1282;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_259 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h103 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_259 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_259 <= _GEN_1283;
      end
    end else begin
      lvtReg_259 <= _GEN_1283;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_260 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h104 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_260 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_260 <= _GEN_1284;
      end
    end else begin
      lvtReg_260 <= _GEN_1284;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_261 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h105 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_261 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_261 <= _GEN_1285;
      end
    end else begin
      lvtReg_261 <= _GEN_1285;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_262 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h106 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_262 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_262 <= _GEN_1286;
      end
    end else begin
      lvtReg_262 <= _GEN_1286;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_263 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h107 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_263 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_263 <= _GEN_1287;
      end
    end else begin
      lvtReg_263 <= _GEN_1287;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_264 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h108 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_264 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_264 <= _GEN_1288;
      end
    end else begin
      lvtReg_264 <= _GEN_1288;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_265 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h109 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_265 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_265 <= _GEN_1289;
      end
    end else begin
      lvtReg_265 <= _GEN_1289;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_266 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_266 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_266 <= _GEN_1290;
      end
    end else begin
      lvtReg_266 <= _GEN_1290;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_267 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_267 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_267 <= _GEN_1291;
      end
    end else begin
      lvtReg_267 <= _GEN_1291;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_268 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_268 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_268 <= _GEN_1292;
      end
    end else begin
      lvtReg_268 <= _GEN_1292;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_269 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_269 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_269 <= _GEN_1293;
      end
    end else begin
      lvtReg_269 <= _GEN_1293;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_270 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_270 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_270 <= _GEN_1294;
      end
    end else begin
      lvtReg_270 <= _GEN_1294;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_271 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h10f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_271 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_271 <= _GEN_1295;
      end
    end else begin
      lvtReg_271 <= _GEN_1295;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_272 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h110 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_272 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_272 <= _GEN_1296;
      end
    end else begin
      lvtReg_272 <= _GEN_1296;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_273 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h111 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_273 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_273 <= _GEN_1297;
      end
    end else begin
      lvtReg_273 <= _GEN_1297;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_274 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h112 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_274 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_274 <= _GEN_1298;
      end
    end else begin
      lvtReg_274 <= _GEN_1298;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_275 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h113 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_275 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_275 <= _GEN_1299;
      end
    end else begin
      lvtReg_275 <= _GEN_1299;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_276 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h114 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_276 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_276 <= _GEN_1300;
      end
    end else begin
      lvtReg_276 <= _GEN_1300;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_277 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h115 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_277 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_277 <= _GEN_1301;
      end
    end else begin
      lvtReg_277 <= _GEN_1301;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_278 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h116 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_278 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_278 <= _GEN_1302;
      end
    end else begin
      lvtReg_278 <= _GEN_1302;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_279 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h117 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_279 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_279 <= _GEN_1303;
      end
    end else begin
      lvtReg_279 <= _GEN_1303;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_280 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h118 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_280 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_280 <= _GEN_1304;
      end
    end else begin
      lvtReg_280 <= _GEN_1304;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_281 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h119 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_281 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_281 <= _GEN_1305;
      end
    end else begin
      lvtReg_281 <= _GEN_1305;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_282 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_282 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_282 <= _GEN_1306;
      end
    end else begin
      lvtReg_282 <= _GEN_1306;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_283 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_283 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_283 <= _GEN_1307;
      end
    end else begin
      lvtReg_283 <= _GEN_1307;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_284 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_284 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_284 <= _GEN_1308;
      end
    end else begin
      lvtReg_284 <= _GEN_1308;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_285 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_285 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_285 <= _GEN_1309;
      end
    end else begin
      lvtReg_285 <= _GEN_1309;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_286 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_286 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_286 <= _GEN_1310;
      end
    end else begin
      lvtReg_286 <= _GEN_1310;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_287 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h11f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_287 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_287 <= _GEN_1311;
      end
    end else begin
      lvtReg_287 <= _GEN_1311;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_288 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h120 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_288 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_288 <= _GEN_1312;
      end
    end else begin
      lvtReg_288 <= _GEN_1312;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_289 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h121 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_289 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_289 <= _GEN_1313;
      end
    end else begin
      lvtReg_289 <= _GEN_1313;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_290 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h122 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_290 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_290 <= _GEN_1314;
      end
    end else begin
      lvtReg_290 <= _GEN_1314;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_291 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h123 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_291 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_291 <= _GEN_1315;
      end
    end else begin
      lvtReg_291 <= _GEN_1315;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_292 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h124 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_292 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_292 <= _GEN_1316;
      end
    end else begin
      lvtReg_292 <= _GEN_1316;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_293 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h125 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_293 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_293 <= _GEN_1317;
      end
    end else begin
      lvtReg_293 <= _GEN_1317;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_294 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h126 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_294 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_294 <= _GEN_1318;
      end
    end else begin
      lvtReg_294 <= _GEN_1318;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_295 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h127 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_295 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_295 <= _GEN_1319;
      end
    end else begin
      lvtReg_295 <= _GEN_1319;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_296 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h128 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_296 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_296 <= _GEN_1320;
      end
    end else begin
      lvtReg_296 <= _GEN_1320;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_297 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h129 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_297 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_297 <= _GEN_1321;
      end
    end else begin
      lvtReg_297 <= _GEN_1321;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_298 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_298 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_298 <= _GEN_1322;
      end
    end else begin
      lvtReg_298 <= _GEN_1322;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_299 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_299 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_299 <= _GEN_1323;
      end
    end else begin
      lvtReg_299 <= _GEN_1323;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_300 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_300 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_300 <= _GEN_1324;
      end
    end else begin
      lvtReg_300 <= _GEN_1324;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_301 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_301 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_301 <= _GEN_1325;
      end
    end else begin
      lvtReg_301 <= _GEN_1325;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_302 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_302 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_302 <= _GEN_1326;
      end
    end else begin
      lvtReg_302 <= _GEN_1326;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_303 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h12f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_303 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_303 <= _GEN_1327;
      end
    end else begin
      lvtReg_303 <= _GEN_1327;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_304 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h130 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_304 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_304 <= _GEN_1328;
      end
    end else begin
      lvtReg_304 <= _GEN_1328;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_305 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h131 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_305 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_305 <= _GEN_1329;
      end
    end else begin
      lvtReg_305 <= _GEN_1329;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_306 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h132 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_306 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_306 <= _GEN_1330;
      end
    end else begin
      lvtReg_306 <= _GEN_1330;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_307 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h133 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_307 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_307 <= _GEN_1331;
      end
    end else begin
      lvtReg_307 <= _GEN_1331;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_308 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h134 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_308 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_308 <= _GEN_1332;
      end
    end else begin
      lvtReg_308 <= _GEN_1332;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_309 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h135 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_309 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_309 <= _GEN_1333;
      end
    end else begin
      lvtReg_309 <= _GEN_1333;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_310 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h136 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_310 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_310 <= _GEN_1334;
      end
    end else begin
      lvtReg_310 <= _GEN_1334;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_311 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h137 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_311 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_311 <= _GEN_1335;
      end
    end else begin
      lvtReg_311 <= _GEN_1335;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_312 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h138 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_312 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_312 <= _GEN_1336;
      end
    end else begin
      lvtReg_312 <= _GEN_1336;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_313 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h139 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_313 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_313 <= _GEN_1337;
      end
    end else begin
      lvtReg_313 <= _GEN_1337;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_314 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_314 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_314 <= _GEN_1338;
      end
    end else begin
      lvtReg_314 <= _GEN_1338;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_315 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_315 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_315 <= _GEN_1339;
      end
    end else begin
      lvtReg_315 <= _GEN_1339;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_316 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_316 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_316 <= _GEN_1340;
      end
    end else begin
      lvtReg_316 <= _GEN_1340;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_317 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_317 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_317 <= _GEN_1341;
      end
    end else begin
      lvtReg_317 <= _GEN_1341;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_318 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_318 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_318 <= _GEN_1342;
      end
    end else begin
      lvtReg_318 <= _GEN_1342;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_319 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h13f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_319 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_319 <= _GEN_1343;
      end
    end else begin
      lvtReg_319 <= _GEN_1343;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_320 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h140 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_320 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_320 <= _GEN_1344;
      end
    end else begin
      lvtReg_320 <= _GEN_1344;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_321 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h141 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_321 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_321 <= _GEN_1345;
      end
    end else begin
      lvtReg_321 <= _GEN_1345;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_322 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h142 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_322 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_322 <= _GEN_1346;
      end
    end else begin
      lvtReg_322 <= _GEN_1346;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_323 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h143 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_323 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_323 <= _GEN_1347;
      end
    end else begin
      lvtReg_323 <= _GEN_1347;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_324 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h144 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_324 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_324 <= _GEN_1348;
      end
    end else begin
      lvtReg_324 <= _GEN_1348;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_325 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h145 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_325 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_325 <= _GEN_1349;
      end
    end else begin
      lvtReg_325 <= _GEN_1349;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_326 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h146 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_326 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_326 <= _GEN_1350;
      end
    end else begin
      lvtReg_326 <= _GEN_1350;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_327 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h147 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_327 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_327 <= _GEN_1351;
      end
    end else begin
      lvtReg_327 <= _GEN_1351;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_328 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h148 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_328 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_328 <= _GEN_1352;
      end
    end else begin
      lvtReg_328 <= _GEN_1352;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_329 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h149 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_329 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_329 <= _GEN_1353;
      end
    end else begin
      lvtReg_329 <= _GEN_1353;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_330 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_330 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_330 <= _GEN_1354;
      end
    end else begin
      lvtReg_330 <= _GEN_1354;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_331 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_331 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_331 <= _GEN_1355;
      end
    end else begin
      lvtReg_331 <= _GEN_1355;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_332 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_332 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_332 <= _GEN_1356;
      end
    end else begin
      lvtReg_332 <= _GEN_1356;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_333 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_333 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_333 <= _GEN_1357;
      end
    end else begin
      lvtReg_333 <= _GEN_1357;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_334 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_334 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_334 <= _GEN_1358;
      end
    end else begin
      lvtReg_334 <= _GEN_1358;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_335 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h14f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_335 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_335 <= _GEN_1359;
      end
    end else begin
      lvtReg_335 <= _GEN_1359;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_336 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h150 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_336 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_336 <= _GEN_1360;
      end
    end else begin
      lvtReg_336 <= _GEN_1360;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_337 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h151 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_337 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_337 <= _GEN_1361;
      end
    end else begin
      lvtReg_337 <= _GEN_1361;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_338 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h152 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_338 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_338 <= _GEN_1362;
      end
    end else begin
      lvtReg_338 <= _GEN_1362;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_339 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h153 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_339 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_339 <= _GEN_1363;
      end
    end else begin
      lvtReg_339 <= _GEN_1363;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_340 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h154 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_340 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_340 <= _GEN_1364;
      end
    end else begin
      lvtReg_340 <= _GEN_1364;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_341 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h155 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_341 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_341 <= _GEN_1365;
      end
    end else begin
      lvtReg_341 <= _GEN_1365;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_342 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h156 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_342 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_342 <= _GEN_1366;
      end
    end else begin
      lvtReg_342 <= _GEN_1366;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_343 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h157 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_343 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_343 <= _GEN_1367;
      end
    end else begin
      lvtReg_343 <= _GEN_1367;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_344 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h158 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_344 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_344 <= _GEN_1368;
      end
    end else begin
      lvtReg_344 <= _GEN_1368;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_345 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h159 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_345 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_345 <= _GEN_1369;
      end
    end else begin
      lvtReg_345 <= _GEN_1369;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_346 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_346 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_346 <= _GEN_1370;
      end
    end else begin
      lvtReg_346 <= _GEN_1370;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_347 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_347 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_347 <= _GEN_1371;
      end
    end else begin
      lvtReg_347 <= _GEN_1371;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_348 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_348 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_348 <= _GEN_1372;
      end
    end else begin
      lvtReg_348 <= _GEN_1372;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_349 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_349 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_349 <= _GEN_1373;
      end
    end else begin
      lvtReg_349 <= _GEN_1373;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_350 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_350 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_350 <= _GEN_1374;
      end
    end else begin
      lvtReg_350 <= _GEN_1374;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_351 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h15f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_351 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_351 <= _GEN_1375;
      end
    end else begin
      lvtReg_351 <= _GEN_1375;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_352 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h160 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_352 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_352 <= _GEN_1376;
      end
    end else begin
      lvtReg_352 <= _GEN_1376;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_353 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h161 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_353 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_353 <= _GEN_1377;
      end
    end else begin
      lvtReg_353 <= _GEN_1377;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_354 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h162 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_354 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_354 <= _GEN_1378;
      end
    end else begin
      lvtReg_354 <= _GEN_1378;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_355 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h163 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_355 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_355 <= _GEN_1379;
      end
    end else begin
      lvtReg_355 <= _GEN_1379;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_356 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h164 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_356 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_356 <= _GEN_1380;
      end
    end else begin
      lvtReg_356 <= _GEN_1380;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_357 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h165 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_357 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_357 <= _GEN_1381;
      end
    end else begin
      lvtReg_357 <= _GEN_1381;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_358 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h166 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_358 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_358 <= _GEN_1382;
      end
    end else begin
      lvtReg_358 <= _GEN_1382;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_359 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h167 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_359 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_359 <= _GEN_1383;
      end
    end else begin
      lvtReg_359 <= _GEN_1383;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_360 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h168 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_360 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_360 <= _GEN_1384;
      end
    end else begin
      lvtReg_360 <= _GEN_1384;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_361 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h169 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_361 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_361 <= _GEN_1385;
      end
    end else begin
      lvtReg_361 <= _GEN_1385;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_362 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_362 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_362 <= _GEN_1386;
      end
    end else begin
      lvtReg_362 <= _GEN_1386;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_363 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_363 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_363 <= _GEN_1387;
      end
    end else begin
      lvtReg_363 <= _GEN_1387;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_364 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_364 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_364 <= _GEN_1388;
      end
    end else begin
      lvtReg_364 <= _GEN_1388;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_365 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_365 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_365 <= _GEN_1389;
      end
    end else begin
      lvtReg_365 <= _GEN_1389;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_366 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_366 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_366 <= _GEN_1390;
      end
    end else begin
      lvtReg_366 <= _GEN_1390;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_367 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h16f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_367 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_367 <= _GEN_1391;
      end
    end else begin
      lvtReg_367 <= _GEN_1391;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_368 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h170 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_368 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_368 <= _GEN_1392;
      end
    end else begin
      lvtReg_368 <= _GEN_1392;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_369 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h171 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_369 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_369 <= _GEN_1393;
      end
    end else begin
      lvtReg_369 <= _GEN_1393;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_370 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h172 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_370 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_370 <= _GEN_1394;
      end
    end else begin
      lvtReg_370 <= _GEN_1394;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_371 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h173 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_371 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_371 <= _GEN_1395;
      end
    end else begin
      lvtReg_371 <= _GEN_1395;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_372 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h174 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_372 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_372 <= _GEN_1396;
      end
    end else begin
      lvtReg_372 <= _GEN_1396;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_373 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h175 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_373 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_373 <= _GEN_1397;
      end
    end else begin
      lvtReg_373 <= _GEN_1397;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_374 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h176 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_374 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_374 <= _GEN_1398;
      end
    end else begin
      lvtReg_374 <= _GEN_1398;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_375 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h177 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_375 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_375 <= _GEN_1399;
      end
    end else begin
      lvtReg_375 <= _GEN_1399;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_376 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h178 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_376 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_376 <= _GEN_1400;
      end
    end else begin
      lvtReg_376 <= _GEN_1400;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_377 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h179 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_377 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_377 <= _GEN_1401;
      end
    end else begin
      lvtReg_377 <= _GEN_1401;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_378 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_378 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_378 <= _GEN_1402;
      end
    end else begin
      lvtReg_378 <= _GEN_1402;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_379 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_379 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_379 <= _GEN_1403;
      end
    end else begin
      lvtReg_379 <= _GEN_1403;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_380 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_380 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_380 <= _GEN_1404;
      end
    end else begin
      lvtReg_380 <= _GEN_1404;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_381 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_381 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_381 <= _GEN_1405;
      end
    end else begin
      lvtReg_381 <= _GEN_1405;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_382 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_382 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_382 <= _GEN_1406;
      end
    end else begin
      lvtReg_382 <= _GEN_1406;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_383 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h17f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_383 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_383 <= _GEN_1407;
      end
    end else begin
      lvtReg_383 <= _GEN_1407;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_384 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h180 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_384 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_384 <= _GEN_1408;
      end
    end else begin
      lvtReg_384 <= _GEN_1408;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_385 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h181 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_385 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_385 <= _GEN_1409;
      end
    end else begin
      lvtReg_385 <= _GEN_1409;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_386 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h182 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_386 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_386 <= _GEN_1410;
      end
    end else begin
      lvtReg_386 <= _GEN_1410;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_387 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h183 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_387 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_387 <= _GEN_1411;
      end
    end else begin
      lvtReg_387 <= _GEN_1411;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_388 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h184 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_388 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_388 <= _GEN_1412;
      end
    end else begin
      lvtReg_388 <= _GEN_1412;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_389 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h185 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_389 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_389 <= _GEN_1413;
      end
    end else begin
      lvtReg_389 <= _GEN_1413;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_390 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h186 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_390 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_390 <= _GEN_1414;
      end
    end else begin
      lvtReg_390 <= _GEN_1414;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_391 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h187 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_391 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_391 <= _GEN_1415;
      end
    end else begin
      lvtReg_391 <= _GEN_1415;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_392 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h188 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_392 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_392 <= _GEN_1416;
      end
    end else begin
      lvtReg_392 <= _GEN_1416;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_393 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h189 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_393 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_393 <= _GEN_1417;
      end
    end else begin
      lvtReg_393 <= _GEN_1417;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_394 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_394 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_394 <= _GEN_1418;
      end
    end else begin
      lvtReg_394 <= _GEN_1418;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_395 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_395 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_395 <= _GEN_1419;
      end
    end else begin
      lvtReg_395 <= _GEN_1419;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_396 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_396 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_396 <= _GEN_1420;
      end
    end else begin
      lvtReg_396 <= _GEN_1420;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_397 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_397 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_397 <= _GEN_1421;
      end
    end else begin
      lvtReg_397 <= _GEN_1421;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_398 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_398 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_398 <= _GEN_1422;
      end
    end else begin
      lvtReg_398 <= _GEN_1422;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_399 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h18f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_399 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_399 <= _GEN_1423;
      end
    end else begin
      lvtReg_399 <= _GEN_1423;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_400 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h190 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_400 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_400 <= _GEN_1424;
      end
    end else begin
      lvtReg_400 <= _GEN_1424;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_401 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h191 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_401 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_401 <= _GEN_1425;
      end
    end else begin
      lvtReg_401 <= _GEN_1425;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_402 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h192 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_402 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_402 <= _GEN_1426;
      end
    end else begin
      lvtReg_402 <= _GEN_1426;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_403 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h193 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_403 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_403 <= _GEN_1427;
      end
    end else begin
      lvtReg_403 <= _GEN_1427;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_404 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h194 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_404 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_404 <= _GEN_1428;
      end
    end else begin
      lvtReg_404 <= _GEN_1428;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_405 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h195 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_405 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_405 <= _GEN_1429;
      end
    end else begin
      lvtReg_405 <= _GEN_1429;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_406 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h196 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_406 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_406 <= _GEN_1430;
      end
    end else begin
      lvtReg_406 <= _GEN_1430;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_407 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h197 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_407 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_407 <= _GEN_1431;
      end
    end else begin
      lvtReg_407 <= _GEN_1431;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_408 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h198 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_408 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_408 <= _GEN_1432;
      end
    end else begin
      lvtReg_408 <= _GEN_1432;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_409 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h199 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_409 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_409 <= _GEN_1433;
      end
    end else begin
      lvtReg_409 <= _GEN_1433;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_410 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_410 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_410 <= _GEN_1434;
      end
    end else begin
      lvtReg_410 <= _GEN_1434;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_411 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_411 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_411 <= _GEN_1435;
      end
    end else begin
      lvtReg_411 <= _GEN_1435;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_412 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_412 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_412 <= _GEN_1436;
      end
    end else begin
      lvtReg_412 <= _GEN_1436;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_413 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_413 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_413 <= _GEN_1437;
      end
    end else begin
      lvtReg_413 <= _GEN_1437;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_414 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_414 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_414 <= _GEN_1438;
      end
    end else begin
      lvtReg_414 <= _GEN_1438;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_415 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h19f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_415 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_415 <= _GEN_1439;
      end
    end else begin
      lvtReg_415 <= _GEN_1439;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_416 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_416 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_416 <= _GEN_1440;
      end
    end else begin
      lvtReg_416 <= _GEN_1440;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_417 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_417 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_417 <= _GEN_1441;
      end
    end else begin
      lvtReg_417 <= _GEN_1441;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_418 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_418 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_418 <= _GEN_1442;
      end
    end else begin
      lvtReg_418 <= _GEN_1442;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_419 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_419 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_419 <= _GEN_1443;
      end
    end else begin
      lvtReg_419 <= _GEN_1443;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_420 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_420 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_420 <= _GEN_1444;
      end
    end else begin
      lvtReg_420 <= _GEN_1444;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_421 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_421 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_421 <= _GEN_1445;
      end
    end else begin
      lvtReg_421 <= _GEN_1445;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_422 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_422 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_422 <= _GEN_1446;
      end
    end else begin
      lvtReg_422 <= _GEN_1446;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_423 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_423 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_423 <= _GEN_1447;
      end
    end else begin
      lvtReg_423 <= _GEN_1447;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_424 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_424 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_424 <= _GEN_1448;
      end
    end else begin
      lvtReg_424 <= _GEN_1448;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_425 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1a9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_425 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_425 <= _GEN_1449;
      end
    end else begin
      lvtReg_425 <= _GEN_1449;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_426 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1aa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_426 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_426 <= _GEN_1450;
      end
    end else begin
      lvtReg_426 <= _GEN_1450;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_427 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ab == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_427 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_427 <= _GEN_1451;
      end
    end else begin
      lvtReg_427 <= _GEN_1451;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_428 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ac == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_428 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_428 <= _GEN_1452;
      end
    end else begin
      lvtReg_428 <= _GEN_1452;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_429 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ad == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_429 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_429 <= _GEN_1453;
      end
    end else begin
      lvtReg_429 <= _GEN_1453;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_430 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ae == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_430 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_430 <= _GEN_1454;
      end
    end else begin
      lvtReg_430 <= _GEN_1454;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_431 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1af == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_431 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_431 <= _GEN_1455;
      end
    end else begin
      lvtReg_431 <= _GEN_1455;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_432 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_432 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_432 <= _GEN_1456;
      end
    end else begin
      lvtReg_432 <= _GEN_1456;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_433 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_433 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_433 <= _GEN_1457;
      end
    end else begin
      lvtReg_433 <= _GEN_1457;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_434 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_434 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_434 <= _GEN_1458;
      end
    end else begin
      lvtReg_434 <= _GEN_1458;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_435 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_435 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_435 <= _GEN_1459;
      end
    end else begin
      lvtReg_435 <= _GEN_1459;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_436 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_436 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_436 <= _GEN_1460;
      end
    end else begin
      lvtReg_436 <= _GEN_1460;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_437 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_437 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_437 <= _GEN_1461;
      end
    end else begin
      lvtReg_437 <= _GEN_1461;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_438 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_438 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_438 <= _GEN_1462;
      end
    end else begin
      lvtReg_438 <= _GEN_1462;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_439 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_439 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_439 <= _GEN_1463;
      end
    end else begin
      lvtReg_439 <= _GEN_1463;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_440 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_440 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_440 <= _GEN_1464;
      end
    end else begin
      lvtReg_440 <= _GEN_1464;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_441 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1b9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_441 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_441 <= _GEN_1465;
      end
    end else begin
      lvtReg_441 <= _GEN_1465;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_442 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ba == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_442 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_442 <= _GEN_1466;
      end
    end else begin
      lvtReg_442 <= _GEN_1466;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_443 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1bb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_443 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_443 <= _GEN_1467;
      end
    end else begin
      lvtReg_443 <= _GEN_1467;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_444 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1bc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_444 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_444 <= _GEN_1468;
      end
    end else begin
      lvtReg_444 <= _GEN_1468;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_445 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1bd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_445 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_445 <= _GEN_1469;
      end
    end else begin
      lvtReg_445 <= _GEN_1469;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_446 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1be == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_446 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_446 <= _GEN_1470;
      end
    end else begin
      lvtReg_446 <= _GEN_1470;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_447 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1bf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_447 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_447 <= _GEN_1471;
      end
    end else begin
      lvtReg_447 <= _GEN_1471;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_448 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_448 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_448 <= _GEN_1472;
      end
    end else begin
      lvtReg_448 <= _GEN_1472;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_449 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_449 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_449 <= _GEN_1473;
      end
    end else begin
      lvtReg_449 <= _GEN_1473;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_450 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_450 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_450 <= _GEN_1474;
      end
    end else begin
      lvtReg_450 <= _GEN_1474;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_451 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_451 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_451 <= _GEN_1475;
      end
    end else begin
      lvtReg_451 <= _GEN_1475;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_452 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_452 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_452 <= _GEN_1476;
      end
    end else begin
      lvtReg_452 <= _GEN_1476;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_453 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_453 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_453 <= _GEN_1477;
      end
    end else begin
      lvtReg_453 <= _GEN_1477;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_454 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_454 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_454 <= _GEN_1478;
      end
    end else begin
      lvtReg_454 <= _GEN_1478;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_455 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_455 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_455 <= _GEN_1479;
      end
    end else begin
      lvtReg_455 <= _GEN_1479;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_456 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_456 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_456 <= _GEN_1480;
      end
    end else begin
      lvtReg_456 <= _GEN_1480;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_457 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1c9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_457 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_457 <= _GEN_1481;
      end
    end else begin
      lvtReg_457 <= _GEN_1481;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_458 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ca == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_458 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_458 <= _GEN_1482;
      end
    end else begin
      lvtReg_458 <= _GEN_1482;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_459 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1cb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_459 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_459 <= _GEN_1483;
      end
    end else begin
      lvtReg_459 <= _GEN_1483;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_460 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1cc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_460 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_460 <= _GEN_1484;
      end
    end else begin
      lvtReg_460 <= _GEN_1484;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_461 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1cd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_461 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_461 <= _GEN_1485;
      end
    end else begin
      lvtReg_461 <= _GEN_1485;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_462 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ce == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_462 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_462 <= _GEN_1486;
      end
    end else begin
      lvtReg_462 <= _GEN_1486;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_463 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1cf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_463 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_463 <= _GEN_1487;
      end
    end else begin
      lvtReg_463 <= _GEN_1487;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_464 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_464 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_464 <= _GEN_1488;
      end
    end else begin
      lvtReg_464 <= _GEN_1488;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_465 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_465 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_465 <= _GEN_1489;
      end
    end else begin
      lvtReg_465 <= _GEN_1489;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_466 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_466 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_466 <= _GEN_1490;
      end
    end else begin
      lvtReg_466 <= _GEN_1490;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_467 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_467 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_467 <= _GEN_1491;
      end
    end else begin
      lvtReg_467 <= _GEN_1491;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_468 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_468 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_468 <= _GEN_1492;
      end
    end else begin
      lvtReg_468 <= _GEN_1492;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_469 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_469 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_469 <= _GEN_1493;
      end
    end else begin
      lvtReg_469 <= _GEN_1493;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_470 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_470 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_470 <= _GEN_1494;
      end
    end else begin
      lvtReg_470 <= _GEN_1494;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_471 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_471 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_471 <= _GEN_1495;
      end
    end else begin
      lvtReg_471 <= _GEN_1495;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_472 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_472 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_472 <= _GEN_1496;
      end
    end else begin
      lvtReg_472 <= _GEN_1496;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_473 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1d9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_473 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_473 <= _GEN_1497;
      end
    end else begin
      lvtReg_473 <= _GEN_1497;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_474 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1da == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_474 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_474 <= _GEN_1498;
      end
    end else begin
      lvtReg_474 <= _GEN_1498;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_475 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1db == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_475 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_475 <= _GEN_1499;
      end
    end else begin
      lvtReg_475 <= _GEN_1499;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_476 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1dc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_476 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_476 <= _GEN_1500;
      end
    end else begin
      lvtReg_476 <= _GEN_1500;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_477 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1dd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_477 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_477 <= _GEN_1501;
      end
    end else begin
      lvtReg_477 <= _GEN_1501;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_478 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1de == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_478 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_478 <= _GEN_1502;
      end
    end else begin
      lvtReg_478 <= _GEN_1502;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_479 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1df == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_479 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_479 <= _GEN_1503;
      end
    end else begin
      lvtReg_479 <= _GEN_1503;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_480 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_480 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_480 <= _GEN_1504;
      end
    end else begin
      lvtReg_480 <= _GEN_1504;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_481 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_481 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_481 <= _GEN_1505;
      end
    end else begin
      lvtReg_481 <= _GEN_1505;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_482 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_482 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_482 <= _GEN_1506;
      end
    end else begin
      lvtReg_482 <= _GEN_1506;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_483 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_483 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_483 <= _GEN_1507;
      end
    end else begin
      lvtReg_483 <= _GEN_1507;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_484 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_484 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_484 <= _GEN_1508;
      end
    end else begin
      lvtReg_484 <= _GEN_1508;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_485 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_485 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_485 <= _GEN_1509;
      end
    end else begin
      lvtReg_485 <= _GEN_1509;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_486 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_486 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_486 <= _GEN_1510;
      end
    end else begin
      lvtReg_486 <= _GEN_1510;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_487 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_487 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_487 <= _GEN_1511;
      end
    end else begin
      lvtReg_487 <= _GEN_1511;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_488 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_488 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_488 <= _GEN_1512;
      end
    end else begin
      lvtReg_488 <= _GEN_1512;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_489 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1e9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_489 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_489 <= _GEN_1513;
      end
    end else begin
      lvtReg_489 <= _GEN_1513;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_490 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ea == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_490 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_490 <= _GEN_1514;
      end
    end else begin
      lvtReg_490 <= _GEN_1514;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_491 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1eb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_491 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_491 <= _GEN_1515;
      end
    end else begin
      lvtReg_491 <= _GEN_1515;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_492 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ec == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_492 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_492 <= _GEN_1516;
      end
    end else begin
      lvtReg_492 <= _GEN_1516;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_493 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ed == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_493 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_493 <= _GEN_1517;
      end
    end else begin
      lvtReg_493 <= _GEN_1517;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_494 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ee == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_494 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_494 <= _GEN_1518;
      end
    end else begin
      lvtReg_494 <= _GEN_1518;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_495 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ef == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_495 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_495 <= _GEN_1519;
      end
    end else begin
      lvtReg_495 <= _GEN_1519;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_496 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_496 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_496 <= _GEN_1520;
      end
    end else begin
      lvtReg_496 <= _GEN_1520;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_497 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_497 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_497 <= _GEN_1521;
      end
    end else begin
      lvtReg_497 <= _GEN_1521;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_498 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_498 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_498 <= _GEN_1522;
      end
    end else begin
      lvtReg_498 <= _GEN_1522;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_499 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_499 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_499 <= _GEN_1523;
      end
    end else begin
      lvtReg_499 <= _GEN_1523;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_500 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_500 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_500 <= _GEN_1524;
      end
    end else begin
      lvtReg_500 <= _GEN_1524;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_501 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_501 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_501 <= _GEN_1525;
      end
    end else begin
      lvtReg_501 <= _GEN_1525;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_502 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_502 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_502 <= _GEN_1526;
      end
    end else begin
      lvtReg_502 <= _GEN_1526;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_503 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_503 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_503 <= _GEN_1527;
      end
    end else begin
      lvtReg_503 <= _GEN_1527;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_504 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_504 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_504 <= _GEN_1528;
      end
    end else begin
      lvtReg_504 <= _GEN_1528;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_505 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1f9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_505 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_505 <= _GEN_1529;
      end
    end else begin
      lvtReg_505 <= _GEN_1529;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_506 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1fa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_506 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_506 <= _GEN_1530;
      end
    end else begin
      lvtReg_506 <= _GEN_1530;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_507 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1fb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_507 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_507 <= _GEN_1531;
      end
    end else begin
      lvtReg_507 <= _GEN_1531;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_508 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1fc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_508 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_508 <= _GEN_1532;
      end
    end else begin
      lvtReg_508 <= _GEN_1532;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_509 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1fd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_509 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_509 <= _GEN_1533;
      end
    end else begin
      lvtReg_509 <= _GEN_1533;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_510 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1fe == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_510 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_510 <= _GEN_1534;
      end
    end else begin
      lvtReg_510 <= _GEN_1534;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_511 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h1ff == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_511 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_511 <= _GEN_1535;
      end
    end else begin
      lvtReg_511 <= _GEN_1535;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_512 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h200 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_512 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_512 <= _GEN_1536;
      end
    end else begin
      lvtReg_512 <= _GEN_1536;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_513 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h201 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_513 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_513 <= _GEN_1537;
      end
    end else begin
      lvtReg_513 <= _GEN_1537;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_514 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h202 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_514 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_514 <= _GEN_1538;
      end
    end else begin
      lvtReg_514 <= _GEN_1538;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_515 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h203 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_515 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_515 <= _GEN_1539;
      end
    end else begin
      lvtReg_515 <= _GEN_1539;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_516 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h204 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_516 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_516 <= _GEN_1540;
      end
    end else begin
      lvtReg_516 <= _GEN_1540;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_517 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h205 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_517 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_517 <= _GEN_1541;
      end
    end else begin
      lvtReg_517 <= _GEN_1541;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_518 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h206 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_518 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_518 <= _GEN_1542;
      end
    end else begin
      lvtReg_518 <= _GEN_1542;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_519 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h207 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_519 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_519 <= _GEN_1543;
      end
    end else begin
      lvtReg_519 <= _GEN_1543;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_520 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h208 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_520 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_520 <= _GEN_1544;
      end
    end else begin
      lvtReg_520 <= _GEN_1544;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_521 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h209 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_521 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_521 <= _GEN_1545;
      end
    end else begin
      lvtReg_521 <= _GEN_1545;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_522 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_522 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_522 <= _GEN_1546;
      end
    end else begin
      lvtReg_522 <= _GEN_1546;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_523 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_523 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_523 <= _GEN_1547;
      end
    end else begin
      lvtReg_523 <= _GEN_1547;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_524 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_524 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_524 <= _GEN_1548;
      end
    end else begin
      lvtReg_524 <= _GEN_1548;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_525 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_525 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_525 <= _GEN_1549;
      end
    end else begin
      lvtReg_525 <= _GEN_1549;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_526 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_526 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_526 <= _GEN_1550;
      end
    end else begin
      lvtReg_526 <= _GEN_1550;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_527 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h20f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_527 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_527 <= _GEN_1551;
      end
    end else begin
      lvtReg_527 <= _GEN_1551;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_528 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h210 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_528 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_528 <= _GEN_1552;
      end
    end else begin
      lvtReg_528 <= _GEN_1552;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_529 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h211 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_529 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_529 <= _GEN_1553;
      end
    end else begin
      lvtReg_529 <= _GEN_1553;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_530 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h212 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_530 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_530 <= _GEN_1554;
      end
    end else begin
      lvtReg_530 <= _GEN_1554;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_531 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h213 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_531 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_531 <= _GEN_1555;
      end
    end else begin
      lvtReg_531 <= _GEN_1555;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_532 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h214 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_532 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_532 <= _GEN_1556;
      end
    end else begin
      lvtReg_532 <= _GEN_1556;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_533 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h215 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_533 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_533 <= _GEN_1557;
      end
    end else begin
      lvtReg_533 <= _GEN_1557;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_534 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h216 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_534 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_534 <= _GEN_1558;
      end
    end else begin
      lvtReg_534 <= _GEN_1558;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_535 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h217 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_535 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_535 <= _GEN_1559;
      end
    end else begin
      lvtReg_535 <= _GEN_1559;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_536 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h218 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_536 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_536 <= _GEN_1560;
      end
    end else begin
      lvtReg_536 <= _GEN_1560;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_537 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h219 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_537 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_537 <= _GEN_1561;
      end
    end else begin
      lvtReg_537 <= _GEN_1561;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_538 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_538 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_538 <= _GEN_1562;
      end
    end else begin
      lvtReg_538 <= _GEN_1562;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_539 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_539 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_539 <= _GEN_1563;
      end
    end else begin
      lvtReg_539 <= _GEN_1563;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_540 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_540 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_540 <= _GEN_1564;
      end
    end else begin
      lvtReg_540 <= _GEN_1564;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_541 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_541 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_541 <= _GEN_1565;
      end
    end else begin
      lvtReg_541 <= _GEN_1565;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_542 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_542 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_542 <= _GEN_1566;
      end
    end else begin
      lvtReg_542 <= _GEN_1566;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_543 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h21f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_543 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_543 <= _GEN_1567;
      end
    end else begin
      lvtReg_543 <= _GEN_1567;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_544 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h220 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_544 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_544 <= _GEN_1568;
      end
    end else begin
      lvtReg_544 <= _GEN_1568;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_545 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h221 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_545 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_545 <= _GEN_1569;
      end
    end else begin
      lvtReg_545 <= _GEN_1569;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_546 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h222 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_546 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_546 <= _GEN_1570;
      end
    end else begin
      lvtReg_546 <= _GEN_1570;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_547 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h223 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_547 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_547 <= _GEN_1571;
      end
    end else begin
      lvtReg_547 <= _GEN_1571;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_548 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h224 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_548 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_548 <= _GEN_1572;
      end
    end else begin
      lvtReg_548 <= _GEN_1572;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_549 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h225 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_549 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_549 <= _GEN_1573;
      end
    end else begin
      lvtReg_549 <= _GEN_1573;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_550 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h226 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_550 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_550 <= _GEN_1574;
      end
    end else begin
      lvtReg_550 <= _GEN_1574;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_551 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h227 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_551 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_551 <= _GEN_1575;
      end
    end else begin
      lvtReg_551 <= _GEN_1575;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_552 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h228 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_552 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_552 <= _GEN_1576;
      end
    end else begin
      lvtReg_552 <= _GEN_1576;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_553 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h229 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_553 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_553 <= _GEN_1577;
      end
    end else begin
      lvtReg_553 <= _GEN_1577;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_554 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_554 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_554 <= _GEN_1578;
      end
    end else begin
      lvtReg_554 <= _GEN_1578;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_555 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_555 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_555 <= _GEN_1579;
      end
    end else begin
      lvtReg_555 <= _GEN_1579;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_556 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_556 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_556 <= _GEN_1580;
      end
    end else begin
      lvtReg_556 <= _GEN_1580;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_557 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_557 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_557 <= _GEN_1581;
      end
    end else begin
      lvtReg_557 <= _GEN_1581;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_558 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_558 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_558 <= _GEN_1582;
      end
    end else begin
      lvtReg_558 <= _GEN_1582;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_559 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h22f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_559 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_559 <= _GEN_1583;
      end
    end else begin
      lvtReg_559 <= _GEN_1583;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_560 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h230 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_560 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_560 <= _GEN_1584;
      end
    end else begin
      lvtReg_560 <= _GEN_1584;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_561 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h231 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_561 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_561 <= _GEN_1585;
      end
    end else begin
      lvtReg_561 <= _GEN_1585;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_562 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h232 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_562 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_562 <= _GEN_1586;
      end
    end else begin
      lvtReg_562 <= _GEN_1586;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_563 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h233 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_563 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_563 <= _GEN_1587;
      end
    end else begin
      lvtReg_563 <= _GEN_1587;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_564 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h234 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_564 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_564 <= _GEN_1588;
      end
    end else begin
      lvtReg_564 <= _GEN_1588;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_565 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h235 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_565 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_565 <= _GEN_1589;
      end
    end else begin
      lvtReg_565 <= _GEN_1589;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_566 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h236 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_566 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_566 <= _GEN_1590;
      end
    end else begin
      lvtReg_566 <= _GEN_1590;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_567 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h237 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_567 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_567 <= _GEN_1591;
      end
    end else begin
      lvtReg_567 <= _GEN_1591;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_568 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h238 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_568 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_568 <= _GEN_1592;
      end
    end else begin
      lvtReg_568 <= _GEN_1592;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_569 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h239 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_569 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_569 <= _GEN_1593;
      end
    end else begin
      lvtReg_569 <= _GEN_1593;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_570 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_570 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_570 <= _GEN_1594;
      end
    end else begin
      lvtReg_570 <= _GEN_1594;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_571 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_571 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_571 <= _GEN_1595;
      end
    end else begin
      lvtReg_571 <= _GEN_1595;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_572 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_572 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_572 <= _GEN_1596;
      end
    end else begin
      lvtReg_572 <= _GEN_1596;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_573 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_573 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_573 <= _GEN_1597;
      end
    end else begin
      lvtReg_573 <= _GEN_1597;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_574 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_574 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_574 <= _GEN_1598;
      end
    end else begin
      lvtReg_574 <= _GEN_1598;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_575 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h23f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_575 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_575 <= _GEN_1599;
      end
    end else begin
      lvtReg_575 <= _GEN_1599;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_576 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h240 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_576 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_576 <= _GEN_1600;
      end
    end else begin
      lvtReg_576 <= _GEN_1600;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_577 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h241 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_577 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_577 <= _GEN_1601;
      end
    end else begin
      lvtReg_577 <= _GEN_1601;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_578 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h242 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_578 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_578 <= _GEN_1602;
      end
    end else begin
      lvtReg_578 <= _GEN_1602;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_579 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h243 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_579 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_579 <= _GEN_1603;
      end
    end else begin
      lvtReg_579 <= _GEN_1603;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_580 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h244 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_580 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_580 <= _GEN_1604;
      end
    end else begin
      lvtReg_580 <= _GEN_1604;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_581 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h245 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_581 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_581 <= _GEN_1605;
      end
    end else begin
      lvtReg_581 <= _GEN_1605;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_582 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h246 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_582 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_582 <= _GEN_1606;
      end
    end else begin
      lvtReg_582 <= _GEN_1606;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_583 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h247 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_583 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_583 <= _GEN_1607;
      end
    end else begin
      lvtReg_583 <= _GEN_1607;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_584 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h248 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_584 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_584 <= _GEN_1608;
      end
    end else begin
      lvtReg_584 <= _GEN_1608;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_585 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h249 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_585 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_585 <= _GEN_1609;
      end
    end else begin
      lvtReg_585 <= _GEN_1609;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_586 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_586 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_586 <= _GEN_1610;
      end
    end else begin
      lvtReg_586 <= _GEN_1610;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_587 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_587 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_587 <= _GEN_1611;
      end
    end else begin
      lvtReg_587 <= _GEN_1611;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_588 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_588 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_588 <= _GEN_1612;
      end
    end else begin
      lvtReg_588 <= _GEN_1612;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_589 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_589 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_589 <= _GEN_1613;
      end
    end else begin
      lvtReg_589 <= _GEN_1613;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_590 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_590 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_590 <= _GEN_1614;
      end
    end else begin
      lvtReg_590 <= _GEN_1614;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_591 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h24f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_591 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_591 <= _GEN_1615;
      end
    end else begin
      lvtReg_591 <= _GEN_1615;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_592 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h250 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_592 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_592 <= _GEN_1616;
      end
    end else begin
      lvtReg_592 <= _GEN_1616;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_593 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h251 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_593 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_593 <= _GEN_1617;
      end
    end else begin
      lvtReg_593 <= _GEN_1617;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_594 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h252 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_594 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_594 <= _GEN_1618;
      end
    end else begin
      lvtReg_594 <= _GEN_1618;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_595 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h253 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_595 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_595 <= _GEN_1619;
      end
    end else begin
      lvtReg_595 <= _GEN_1619;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_596 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h254 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_596 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_596 <= _GEN_1620;
      end
    end else begin
      lvtReg_596 <= _GEN_1620;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_597 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h255 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_597 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_597 <= _GEN_1621;
      end
    end else begin
      lvtReg_597 <= _GEN_1621;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_598 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h256 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_598 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_598 <= _GEN_1622;
      end
    end else begin
      lvtReg_598 <= _GEN_1622;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_599 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h257 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_599 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_599 <= _GEN_1623;
      end
    end else begin
      lvtReg_599 <= _GEN_1623;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_600 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h258 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_600 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_600 <= _GEN_1624;
      end
    end else begin
      lvtReg_600 <= _GEN_1624;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_601 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h259 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_601 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_601 <= _GEN_1625;
      end
    end else begin
      lvtReg_601 <= _GEN_1625;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_602 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_602 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_602 <= _GEN_1626;
      end
    end else begin
      lvtReg_602 <= _GEN_1626;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_603 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_603 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_603 <= _GEN_1627;
      end
    end else begin
      lvtReg_603 <= _GEN_1627;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_604 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_604 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_604 <= _GEN_1628;
      end
    end else begin
      lvtReg_604 <= _GEN_1628;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_605 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_605 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_605 <= _GEN_1629;
      end
    end else begin
      lvtReg_605 <= _GEN_1629;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_606 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_606 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_606 <= _GEN_1630;
      end
    end else begin
      lvtReg_606 <= _GEN_1630;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_607 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h25f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_607 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_607 <= _GEN_1631;
      end
    end else begin
      lvtReg_607 <= _GEN_1631;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_608 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h260 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_608 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_608 <= _GEN_1632;
      end
    end else begin
      lvtReg_608 <= _GEN_1632;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_609 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h261 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_609 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_609 <= _GEN_1633;
      end
    end else begin
      lvtReg_609 <= _GEN_1633;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_610 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h262 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_610 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_610 <= _GEN_1634;
      end
    end else begin
      lvtReg_610 <= _GEN_1634;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_611 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h263 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_611 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_611 <= _GEN_1635;
      end
    end else begin
      lvtReg_611 <= _GEN_1635;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_612 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h264 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_612 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_612 <= _GEN_1636;
      end
    end else begin
      lvtReg_612 <= _GEN_1636;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_613 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h265 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_613 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_613 <= _GEN_1637;
      end
    end else begin
      lvtReg_613 <= _GEN_1637;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_614 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h266 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_614 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_614 <= _GEN_1638;
      end
    end else begin
      lvtReg_614 <= _GEN_1638;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_615 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h267 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_615 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_615 <= _GEN_1639;
      end
    end else begin
      lvtReg_615 <= _GEN_1639;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_616 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h268 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_616 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_616 <= _GEN_1640;
      end
    end else begin
      lvtReg_616 <= _GEN_1640;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_617 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h269 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_617 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_617 <= _GEN_1641;
      end
    end else begin
      lvtReg_617 <= _GEN_1641;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_618 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_618 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_618 <= _GEN_1642;
      end
    end else begin
      lvtReg_618 <= _GEN_1642;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_619 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_619 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_619 <= _GEN_1643;
      end
    end else begin
      lvtReg_619 <= _GEN_1643;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_620 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_620 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_620 <= _GEN_1644;
      end
    end else begin
      lvtReg_620 <= _GEN_1644;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_621 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_621 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_621 <= _GEN_1645;
      end
    end else begin
      lvtReg_621 <= _GEN_1645;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_622 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_622 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_622 <= _GEN_1646;
      end
    end else begin
      lvtReg_622 <= _GEN_1646;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_623 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h26f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_623 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_623 <= _GEN_1647;
      end
    end else begin
      lvtReg_623 <= _GEN_1647;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_624 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h270 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_624 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_624 <= _GEN_1648;
      end
    end else begin
      lvtReg_624 <= _GEN_1648;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_625 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h271 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_625 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_625 <= _GEN_1649;
      end
    end else begin
      lvtReg_625 <= _GEN_1649;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_626 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h272 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_626 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_626 <= _GEN_1650;
      end
    end else begin
      lvtReg_626 <= _GEN_1650;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_627 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h273 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_627 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_627 <= _GEN_1651;
      end
    end else begin
      lvtReg_627 <= _GEN_1651;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_628 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h274 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_628 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_628 <= _GEN_1652;
      end
    end else begin
      lvtReg_628 <= _GEN_1652;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_629 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h275 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_629 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_629 <= _GEN_1653;
      end
    end else begin
      lvtReg_629 <= _GEN_1653;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_630 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h276 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_630 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_630 <= _GEN_1654;
      end
    end else begin
      lvtReg_630 <= _GEN_1654;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_631 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h277 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_631 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_631 <= _GEN_1655;
      end
    end else begin
      lvtReg_631 <= _GEN_1655;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_632 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h278 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_632 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_632 <= _GEN_1656;
      end
    end else begin
      lvtReg_632 <= _GEN_1656;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_633 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h279 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_633 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_633 <= _GEN_1657;
      end
    end else begin
      lvtReg_633 <= _GEN_1657;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_634 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_634 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_634 <= _GEN_1658;
      end
    end else begin
      lvtReg_634 <= _GEN_1658;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_635 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_635 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_635 <= _GEN_1659;
      end
    end else begin
      lvtReg_635 <= _GEN_1659;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_636 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_636 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_636 <= _GEN_1660;
      end
    end else begin
      lvtReg_636 <= _GEN_1660;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_637 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_637 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_637 <= _GEN_1661;
      end
    end else begin
      lvtReg_637 <= _GEN_1661;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_638 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_638 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_638 <= _GEN_1662;
      end
    end else begin
      lvtReg_638 <= _GEN_1662;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_639 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h27f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_639 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_639 <= _GEN_1663;
      end
    end else begin
      lvtReg_639 <= _GEN_1663;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_640 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h280 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_640 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_640 <= _GEN_1664;
      end
    end else begin
      lvtReg_640 <= _GEN_1664;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_641 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h281 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_641 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_641 <= _GEN_1665;
      end
    end else begin
      lvtReg_641 <= _GEN_1665;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_642 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h282 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_642 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_642 <= _GEN_1666;
      end
    end else begin
      lvtReg_642 <= _GEN_1666;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_643 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h283 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_643 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_643 <= _GEN_1667;
      end
    end else begin
      lvtReg_643 <= _GEN_1667;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_644 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h284 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_644 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_644 <= _GEN_1668;
      end
    end else begin
      lvtReg_644 <= _GEN_1668;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_645 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h285 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_645 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_645 <= _GEN_1669;
      end
    end else begin
      lvtReg_645 <= _GEN_1669;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_646 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h286 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_646 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_646 <= _GEN_1670;
      end
    end else begin
      lvtReg_646 <= _GEN_1670;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_647 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h287 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_647 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_647 <= _GEN_1671;
      end
    end else begin
      lvtReg_647 <= _GEN_1671;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_648 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h288 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_648 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_648 <= _GEN_1672;
      end
    end else begin
      lvtReg_648 <= _GEN_1672;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_649 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h289 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_649 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_649 <= _GEN_1673;
      end
    end else begin
      lvtReg_649 <= _GEN_1673;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_650 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_650 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_650 <= _GEN_1674;
      end
    end else begin
      lvtReg_650 <= _GEN_1674;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_651 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_651 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_651 <= _GEN_1675;
      end
    end else begin
      lvtReg_651 <= _GEN_1675;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_652 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_652 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_652 <= _GEN_1676;
      end
    end else begin
      lvtReg_652 <= _GEN_1676;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_653 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_653 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_653 <= _GEN_1677;
      end
    end else begin
      lvtReg_653 <= _GEN_1677;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_654 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_654 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_654 <= _GEN_1678;
      end
    end else begin
      lvtReg_654 <= _GEN_1678;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_655 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h28f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_655 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_655 <= _GEN_1679;
      end
    end else begin
      lvtReg_655 <= _GEN_1679;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_656 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h290 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_656 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_656 <= _GEN_1680;
      end
    end else begin
      lvtReg_656 <= _GEN_1680;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_657 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h291 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_657 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_657 <= _GEN_1681;
      end
    end else begin
      lvtReg_657 <= _GEN_1681;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_658 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h292 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_658 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_658 <= _GEN_1682;
      end
    end else begin
      lvtReg_658 <= _GEN_1682;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_659 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h293 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_659 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_659 <= _GEN_1683;
      end
    end else begin
      lvtReg_659 <= _GEN_1683;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_660 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h294 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_660 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_660 <= _GEN_1684;
      end
    end else begin
      lvtReg_660 <= _GEN_1684;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_661 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h295 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_661 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_661 <= _GEN_1685;
      end
    end else begin
      lvtReg_661 <= _GEN_1685;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_662 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h296 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_662 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_662 <= _GEN_1686;
      end
    end else begin
      lvtReg_662 <= _GEN_1686;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_663 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h297 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_663 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_663 <= _GEN_1687;
      end
    end else begin
      lvtReg_663 <= _GEN_1687;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_664 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h298 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_664 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_664 <= _GEN_1688;
      end
    end else begin
      lvtReg_664 <= _GEN_1688;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_665 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h299 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_665 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_665 <= _GEN_1689;
      end
    end else begin
      lvtReg_665 <= _GEN_1689;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_666 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_666 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_666 <= _GEN_1690;
      end
    end else begin
      lvtReg_666 <= _GEN_1690;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_667 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_667 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_667 <= _GEN_1691;
      end
    end else begin
      lvtReg_667 <= _GEN_1691;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_668 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_668 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_668 <= _GEN_1692;
      end
    end else begin
      lvtReg_668 <= _GEN_1692;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_669 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_669 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_669 <= _GEN_1693;
      end
    end else begin
      lvtReg_669 <= _GEN_1693;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_670 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_670 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_670 <= _GEN_1694;
      end
    end else begin
      lvtReg_670 <= _GEN_1694;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_671 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h29f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_671 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_671 <= _GEN_1695;
      end
    end else begin
      lvtReg_671 <= _GEN_1695;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_672 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_672 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_672 <= _GEN_1696;
      end
    end else begin
      lvtReg_672 <= _GEN_1696;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_673 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_673 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_673 <= _GEN_1697;
      end
    end else begin
      lvtReg_673 <= _GEN_1697;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_674 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_674 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_674 <= _GEN_1698;
      end
    end else begin
      lvtReg_674 <= _GEN_1698;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_675 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_675 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_675 <= _GEN_1699;
      end
    end else begin
      lvtReg_675 <= _GEN_1699;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_676 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_676 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_676 <= _GEN_1700;
      end
    end else begin
      lvtReg_676 <= _GEN_1700;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_677 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_677 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_677 <= _GEN_1701;
      end
    end else begin
      lvtReg_677 <= _GEN_1701;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_678 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_678 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_678 <= _GEN_1702;
      end
    end else begin
      lvtReg_678 <= _GEN_1702;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_679 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_679 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_679 <= _GEN_1703;
      end
    end else begin
      lvtReg_679 <= _GEN_1703;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_680 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_680 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_680 <= _GEN_1704;
      end
    end else begin
      lvtReg_680 <= _GEN_1704;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_681 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2a9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_681 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_681 <= _GEN_1705;
      end
    end else begin
      lvtReg_681 <= _GEN_1705;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_682 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2aa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_682 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_682 <= _GEN_1706;
      end
    end else begin
      lvtReg_682 <= _GEN_1706;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_683 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ab == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_683 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_683 <= _GEN_1707;
      end
    end else begin
      lvtReg_683 <= _GEN_1707;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_684 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ac == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_684 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_684 <= _GEN_1708;
      end
    end else begin
      lvtReg_684 <= _GEN_1708;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_685 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ad == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_685 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_685 <= _GEN_1709;
      end
    end else begin
      lvtReg_685 <= _GEN_1709;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_686 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ae == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_686 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_686 <= _GEN_1710;
      end
    end else begin
      lvtReg_686 <= _GEN_1710;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_687 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2af == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_687 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_687 <= _GEN_1711;
      end
    end else begin
      lvtReg_687 <= _GEN_1711;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_688 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_688 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_688 <= _GEN_1712;
      end
    end else begin
      lvtReg_688 <= _GEN_1712;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_689 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_689 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_689 <= _GEN_1713;
      end
    end else begin
      lvtReg_689 <= _GEN_1713;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_690 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_690 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_690 <= _GEN_1714;
      end
    end else begin
      lvtReg_690 <= _GEN_1714;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_691 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_691 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_691 <= _GEN_1715;
      end
    end else begin
      lvtReg_691 <= _GEN_1715;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_692 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_692 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_692 <= _GEN_1716;
      end
    end else begin
      lvtReg_692 <= _GEN_1716;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_693 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_693 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_693 <= _GEN_1717;
      end
    end else begin
      lvtReg_693 <= _GEN_1717;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_694 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_694 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_694 <= _GEN_1718;
      end
    end else begin
      lvtReg_694 <= _GEN_1718;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_695 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_695 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_695 <= _GEN_1719;
      end
    end else begin
      lvtReg_695 <= _GEN_1719;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_696 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_696 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_696 <= _GEN_1720;
      end
    end else begin
      lvtReg_696 <= _GEN_1720;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_697 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2b9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_697 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_697 <= _GEN_1721;
      end
    end else begin
      lvtReg_697 <= _GEN_1721;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_698 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ba == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_698 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_698 <= _GEN_1722;
      end
    end else begin
      lvtReg_698 <= _GEN_1722;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_699 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2bb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_699 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_699 <= _GEN_1723;
      end
    end else begin
      lvtReg_699 <= _GEN_1723;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_700 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2bc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_700 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_700 <= _GEN_1724;
      end
    end else begin
      lvtReg_700 <= _GEN_1724;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_701 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2bd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_701 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_701 <= _GEN_1725;
      end
    end else begin
      lvtReg_701 <= _GEN_1725;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_702 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2be == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_702 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_702 <= _GEN_1726;
      end
    end else begin
      lvtReg_702 <= _GEN_1726;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_703 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2bf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_703 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_703 <= _GEN_1727;
      end
    end else begin
      lvtReg_703 <= _GEN_1727;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_704 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_704 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_704 <= _GEN_1728;
      end
    end else begin
      lvtReg_704 <= _GEN_1728;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_705 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_705 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_705 <= _GEN_1729;
      end
    end else begin
      lvtReg_705 <= _GEN_1729;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_706 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_706 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_706 <= _GEN_1730;
      end
    end else begin
      lvtReg_706 <= _GEN_1730;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_707 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_707 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_707 <= _GEN_1731;
      end
    end else begin
      lvtReg_707 <= _GEN_1731;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_708 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_708 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_708 <= _GEN_1732;
      end
    end else begin
      lvtReg_708 <= _GEN_1732;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_709 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_709 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_709 <= _GEN_1733;
      end
    end else begin
      lvtReg_709 <= _GEN_1733;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_710 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_710 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_710 <= _GEN_1734;
      end
    end else begin
      lvtReg_710 <= _GEN_1734;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_711 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_711 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_711 <= _GEN_1735;
      end
    end else begin
      lvtReg_711 <= _GEN_1735;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_712 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_712 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_712 <= _GEN_1736;
      end
    end else begin
      lvtReg_712 <= _GEN_1736;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_713 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2c9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_713 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_713 <= _GEN_1737;
      end
    end else begin
      lvtReg_713 <= _GEN_1737;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_714 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ca == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_714 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_714 <= _GEN_1738;
      end
    end else begin
      lvtReg_714 <= _GEN_1738;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_715 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2cb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_715 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_715 <= _GEN_1739;
      end
    end else begin
      lvtReg_715 <= _GEN_1739;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_716 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2cc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_716 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_716 <= _GEN_1740;
      end
    end else begin
      lvtReg_716 <= _GEN_1740;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_717 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2cd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_717 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_717 <= _GEN_1741;
      end
    end else begin
      lvtReg_717 <= _GEN_1741;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_718 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ce == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_718 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_718 <= _GEN_1742;
      end
    end else begin
      lvtReg_718 <= _GEN_1742;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_719 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2cf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_719 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_719 <= _GEN_1743;
      end
    end else begin
      lvtReg_719 <= _GEN_1743;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_720 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_720 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_720 <= _GEN_1744;
      end
    end else begin
      lvtReg_720 <= _GEN_1744;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_721 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_721 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_721 <= _GEN_1745;
      end
    end else begin
      lvtReg_721 <= _GEN_1745;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_722 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_722 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_722 <= _GEN_1746;
      end
    end else begin
      lvtReg_722 <= _GEN_1746;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_723 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_723 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_723 <= _GEN_1747;
      end
    end else begin
      lvtReg_723 <= _GEN_1747;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_724 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_724 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_724 <= _GEN_1748;
      end
    end else begin
      lvtReg_724 <= _GEN_1748;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_725 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_725 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_725 <= _GEN_1749;
      end
    end else begin
      lvtReg_725 <= _GEN_1749;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_726 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_726 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_726 <= _GEN_1750;
      end
    end else begin
      lvtReg_726 <= _GEN_1750;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_727 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_727 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_727 <= _GEN_1751;
      end
    end else begin
      lvtReg_727 <= _GEN_1751;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_728 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_728 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_728 <= _GEN_1752;
      end
    end else begin
      lvtReg_728 <= _GEN_1752;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_729 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2d9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_729 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_729 <= _GEN_1753;
      end
    end else begin
      lvtReg_729 <= _GEN_1753;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_730 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2da == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_730 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_730 <= _GEN_1754;
      end
    end else begin
      lvtReg_730 <= _GEN_1754;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_731 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2db == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_731 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_731 <= _GEN_1755;
      end
    end else begin
      lvtReg_731 <= _GEN_1755;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_732 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2dc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_732 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_732 <= _GEN_1756;
      end
    end else begin
      lvtReg_732 <= _GEN_1756;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_733 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2dd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_733 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_733 <= _GEN_1757;
      end
    end else begin
      lvtReg_733 <= _GEN_1757;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_734 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2de == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_734 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_734 <= _GEN_1758;
      end
    end else begin
      lvtReg_734 <= _GEN_1758;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_735 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2df == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_735 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_735 <= _GEN_1759;
      end
    end else begin
      lvtReg_735 <= _GEN_1759;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_736 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_736 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_736 <= _GEN_1760;
      end
    end else begin
      lvtReg_736 <= _GEN_1760;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_737 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_737 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_737 <= _GEN_1761;
      end
    end else begin
      lvtReg_737 <= _GEN_1761;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_738 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_738 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_738 <= _GEN_1762;
      end
    end else begin
      lvtReg_738 <= _GEN_1762;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_739 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_739 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_739 <= _GEN_1763;
      end
    end else begin
      lvtReg_739 <= _GEN_1763;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_740 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_740 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_740 <= _GEN_1764;
      end
    end else begin
      lvtReg_740 <= _GEN_1764;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_741 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_741 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_741 <= _GEN_1765;
      end
    end else begin
      lvtReg_741 <= _GEN_1765;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_742 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_742 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_742 <= _GEN_1766;
      end
    end else begin
      lvtReg_742 <= _GEN_1766;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_743 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_743 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_743 <= _GEN_1767;
      end
    end else begin
      lvtReg_743 <= _GEN_1767;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_744 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_744 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_744 <= _GEN_1768;
      end
    end else begin
      lvtReg_744 <= _GEN_1768;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_745 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2e9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_745 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_745 <= _GEN_1769;
      end
    end else begin
      lvtReg_745 <= _GEN_1769;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_746 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ea == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_746 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_746 <= _GEN_1770;
      end
    end else begin
      lvtReg_746 <= _GEN_1770;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_747 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2eb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_747 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_747 <= _GEN_1771;
      end
    end else begin
      lvtReg_747 <= _GEN_1771;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_748 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ec == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_748 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_748 <= _GEN_1772;
      end
    end else begin
      lvtReg_748 <= _GEN_1772;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_749 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ed == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_749 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_749 <= _GEN_1773;
      end
    end else begin
      lvtReg_749 <= _GEN_1773;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_750 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ee == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_750 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_750 <= _GEN_1774;
      end
    end else begin
      lvtReg_750 <= _GEN_1774;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_751 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ef == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_751 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_751 <= _GEN_1775;
      end
    end else begin
      lvtReg_751 <= _GEN_1775;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_752 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_752 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_752 <= _GEN_1776;
      end
    end else begin
      lvtReg_752 <= _GEN_1776;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_753 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_753 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_753 <= _GEN_1777;
      end
    end else begin
      lvtReg_753 <= _GEN_1777;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_754 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_754 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_754 <= _GEN_1778;
      end
    end else begin
      lvtReg_754 <= _GEN_1778;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_755 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_755 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_755 <= _GEN_1779;
      end
    end else begin
      lvtReg_755 <= _GEN_1779;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_756 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_756 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_756 <= _GEN_1780;
      end
    end else begin
      lvtReg_756 <= _GEN_1780;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_757 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_757 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_757 <= _GEN_1781;
      end
    end else begin
      lvtReg_757 <= _GEN_1781;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_758 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_758 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_758 <= _GEN_1782;
      end
    end else begin
      lvtReg_758 <= _GEN_1782;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_759 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_759 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_759 <= _GEN_1783;
      end
    end else begin
      lvtReg_759 <= _GEN_1783;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_760 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_760 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_760 <= _GEN_1784;
      end
    end else begin
      lvtReg_760 <= _GEN_1784;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_761 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2f9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_761 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_761 <= _GEN_1785;
      end
    end else begin
      lvtReg_761 <= _GEN_1785;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_762 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2fa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_762 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_762 <= _GEN_1786;
      end
    end else begin
      lvtReg_762 <= _GEN_1786;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_763 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2fb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_763 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_763 <= _GEN_1787;
      end
    end else begin
      lvtReg_763 <= _GEN_1787;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_764 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2fc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_764 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_764 <= _GEN_1788;
      end
    end else begin
      lvtReg_764 <= _GEN_1788;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_765 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2fd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_765 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_765 <= _GEN_1789;
      end
    end else begin
      lvtReg_765 <= _GEN_1789;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_766 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2fe == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_766 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_766 <= _GEN_1790;
      end
    end else begin
      lvtReg_766 <= _GEN_1790;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_767 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h2ff == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_767 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_767 <= _GEN_1791;
      end
    end else begin
      lvtReg_767 <= _GEN_1791;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_768 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h300 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_768 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_768 <= _GEN_1792;
      end
    end else begin
      lvtReg_768 <= _GEN_1792;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_769 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h301 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_769 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_769 <= _GEN_1793;
      end
    end else begin
      lvtReg_769 <= _GEN_1793;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_770 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h302 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_770 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_770 <= _GEN_1794;
      end
    end else begin
      lvtReg_770 <= _GEN_1794;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_771 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h303 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_771 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_771 <= _GEN_1795;
      end
    end else begin
      lvtReg_771 <= _GEN_1795;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_772 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h304 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_772 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_772 <= _GEN_1796;
      end
    end else begin
      lvtReg_772 <= _GEN_1796;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_773 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h305 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_773 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_773 <= _GEN_1797;
      end
    end else begin
      lvtReg_773 <= _GEN_1797;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_774 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h306 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_774 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_774 <= _GEN_1798;
      end
    end else begin
      lvtReg_774 <= _GEN_1798;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_775 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h307 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_775 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_775 <= _GEN_1799;
      end
    end else begin
      lvtReg_775 <= _GEN_1799;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_776 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h308 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_776 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_776 <= _GEN_1800;
      end
    end else begin
      lvtReg_776 <= _GEN_1800;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_777 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h309 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_777 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_777 <= _GEN_1801;
      end
    end else begin
      lvtReg_777 <= _GEN_1801;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_778 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_778 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_778 <= _GEN_1802;
      end
    end else begin
      lvtReg_778 <= _GEN_1802;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_779 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_779 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_779 <= _GEN_1803;
      end
    end else begin
      lvtReg_779 <= _GEN_1803;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_780 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_780 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_780 <= _GEN_1804;
      end
    end else begin
      lvtReg_780 <= _GEN_1804;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_781 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_781 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_781 <= _GEN_1805;
      end
    end else begin
      lvtReg_781 <= _GEN_1805;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_782 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_782 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_782 <= _GEN_1806;
      end
    end else begin
      lvtReg_782 <= _GEN_1806;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_783 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h30f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_783 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_783 <= _GEN_1807;
      end
    end else begin
      lvtReg_783 <= _GEN_1807;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_784 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h310 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_784 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_784 <= _GEN_1808;
      end
    end else begin
      lvtReg_784 <= _GEN_1808;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_785 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h311 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_785 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_785 <= _GEN_1809;
      end
    end else begin
      lvtReg_785 <= _GEN_1809;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_786 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h312 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_786 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_786 <= _GEN_1810;
      end
    end else begin
      lvtReg_786 <= _GEN_1810;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_787 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h313 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_787 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_787 <= _GEN_1811;
      end
    end else begin
      lvtReg_787 <= _GEN_1811;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_788 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h314 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_788 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_788 <= _GEN_1812;
      end
    end else begin
      lvtReg_788 <= _GEN_1812;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_789 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h315 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_789 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_789 <= _GEN_1813;
      end
    end else begin
      lvtReg_789 <= _GEN_1813;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_790 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h316 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_790 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_790 <= _GEN_1814;
      end
    end else begin
      lvtReg_790 <= _GEN_1814;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_791 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h317 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_791 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_791 <= _GEN_1815;
      end
    end else begin
      lvtReg_791 <= _GEN_1815;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_792 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h318 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_792 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_792 <= _GEN_1816;
      end
    end else begin
      lvtReg_792 <= _GEN_1816;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_793 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h319 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_793 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_793 <= _GEN_1817;
      end
    end else begin
      lvtReg_793 <= _GEN_1817;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_794 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_794 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_794 <= _GEN_1818;
      end
    end else begin
      lvtReg_794 <= _GEN_1818;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_795 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_795 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_795 <= _GEN_1819;
      end
    end else begin
      lvtReg_795 <= _GEN_1819;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_796 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_796 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_796 <= _GEN_1820;
      end
    end else begin
      lvtReg_796 <= _GEN_1820;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_797 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_797 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_797 <= _GEN_1821;
      end
    end else begin
      lvtReg_797 <= _GEN_1821;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_798 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_798 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_798 <= _GEN_1822;
      end
    end else begin
      lvtReg_798 <= _GEN_1822;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_799 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h31f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_799 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_799 <= _GEN_1823;
      end
    end else begin
      lvtReg_799 <= _GEN_1823;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_800 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h320 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_800 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_800 <= _GEN_1824;
      end
    end else begin
      lvtReg_800 <= _GEN_1824;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_801 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h321 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_801 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_801 <= _GEN_1825;
      end
    end else begin
      lvtReg_801 <= _GEN_1825;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_802 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h322 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_802 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_802 <= _GEN_1826;
      end
    end else begin
      lvtReg_802 <= _GEN_1826;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_803 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h323 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_803 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_803 <= _GEN_1827;
      end
    end else begin
      lvtReg_803 <= _GEN_1827;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_804 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h324 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_804 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_804 <= _GEN_1828;
      end
    end else begin
      lvtReg_804 <= _GEN_1828;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_805 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h325 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_805 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_805 <= _GEN_1829;
      end
    end else begin
      lvtReg_805 <= _GEN_1829;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_806 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h326 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_806 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_806 <= _GEN_1830;
      end
    end else begin
      lvtReg_806 <= _GEN_1830;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_807 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h327 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_807 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_807 <= _GEN_1831;
      end
    end else begin
      lvtReg_807 <= _GEN_1831;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_808 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h328 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_808 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_808 <= _GEN_1832;
      end
    end else begin
      lvtReg_808 <= _GEN_1832;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_809 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h329 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_809 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_809 <= _GEN_1833;
      end
    end else begin
      lvtReg_809 <= _GEN_1833;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_810 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_810 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_810 <= _GEN_1834;
      end
    end else begin
      lvtReg_810 <= _GEN_1834;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_811 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_811 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_811 <= _GEN_1835;
      end
    end else begin
      lvtReg_811 <= _GEN_1835;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_812 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_812 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_812 <= _GEN_1836;
      end
    end else begin
      lvtReg_812 <= _GEN_1836;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_813 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_813 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_813 <= _GEN_1837;
      end
    end else begin
      lvtReg_813 <= _GEN_1837;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_814 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_814 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_814 <= _GEN_1838;
      end
    end else begin
      lvtReg_814 <= _GEN_1838;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_815 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h32f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_815 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_815 <= _GEN_1839;
      end
    end else begin
      lvtReg_815 <= _GEN_1839;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_816 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h330 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_816 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_816 <= _GEN_1840;
      end
    end else begin
      lvtReg_816 <= _GEN_1840;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_817 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h331 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_817 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_817 <= _GEN_1841;
      end
    end else begin
      lvtReg_817 <= _GEN_1841;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_818 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h332 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_818 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_818 <= _GEN_1842;
      end
    end else begin
      lvtReg_818 <= _GEN_1842;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_819 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h333 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_819 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_819 <= _GEN_1843;
      end
    end else begin
      lvtReg_819 <= _GEN_1843;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_820 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h334 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_820 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_820 <= _GEN_1844;
      end
    end else begin
      lvtReg_820 <= _GEN_1844;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_821 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h335 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_821 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_821 <= _GEN_1845;
      end
    end else begin
      lvtReg_821 <= _GEN_1845;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_822 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h336 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_822 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_822 <= _GEN_1846;
      end
    end else begin
      lvtReg_822 <= _GEN_1846;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_823 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h337 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_823 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_823 <= _GEN_1847;
      end
    end else begin
      lvtReg_823 <= _GEN_1847;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_824 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h338 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_824 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_824 <= _GEN_1848;
      end
    end else begin
      lvtReg_824 <= _GEN_1848;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_825 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h339 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_825 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_825 <= _GEN_1849;
      end
    end else begin
      lvtReg_825 <= _GEN_1849;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_826 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_826 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_826 <= _GEN_1850;
      end
    end else begin
      lvtReg_826 <= _GEN_1850;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_827 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_827 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_827 <= _GEN_1851;
      end
    end else begin
      lvtReg_827 <= _GEN_1851;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_828 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_828 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_828 <= _GEN_1852;
      end
    end else begin
      lvtReg_828 <= _GEN_1852;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_829 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_829 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_829 <= _GEN_1853;
      end
    end else begin
      lvtReg_829 <= _GEN_1853;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_830 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_830 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_830 <= _GEN_1854;
      end
    end else begin
      lvtReg_830 <= _GEN_1854;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_831 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h33f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_831 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_831 <= _GEN_1855;
      end
    end else begin
      lvtReg_831 <= _GEN_1855;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_832 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h340 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_832 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_832 <= _GEN_1856;
      end
    end else begin
      lvtReg_832 <= _GEN_1856;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_833 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h341 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_833 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_833 <= _GEN_1857;
      end
    end else begin
      lvtReg_833 <= _GEN_1857;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_834 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h342 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_834 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_834 <= _GEN_1858;
      end
    end else begin
      lvtReg_834 <= _GEN_1858;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_835 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h343 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_835 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_835 <= _GEN_1859;
      end
    end else begin
      lvtReg_835 <= _GEN_1859;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_836 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h344 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_836 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_836 <= _GEN_1860;
      end
    end else begin
      lvtReg_836 <= _GEN_1860;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_837 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h345 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_837 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_837 <= _GEN_1861;
      end
    end else begin
      lvtReg_837 <= _GEN_1861;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_838 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h346 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_838 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_838 <= _GEN_1862;
      end
    end else begin
      lvtReg_838 <= _GEN_1862;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_839 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h347 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_839 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_839 <= _GEN_1863;
      end
    end else begin
      lvtReg_839 <= _GEN_1863;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_840 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h348 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_840 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_840 <= _GEN_1864;
      end
    end else begin
      lvtReg_840 <= _GEN_1864;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_841 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h349 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_841 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_841 <= _GEN_1865;
      end
    end else begin
      lvtReg_841 <= _GEN_1865;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_842 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_842 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_842 <= _GEN_1866;
      end
    end else begin
      lvtReg_842 <= _GEN_1866;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_843 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_843 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_843 <= _GEN_1867;
      end
    end else begin
      lvtReg_843 <= _GEN_1867;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_844 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_844 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_844 <= _GEN_1868;
      end
    end else begin
      lvtReg_844 <= _GEN_1868;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_845 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_845 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_845 <= _GEN_1869;
      end
    end else begin
      lvtReg_845 <= _GEN_1869;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_846 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_846 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_846 <= _GEN_1870;
      end
    end else begin
      lvtReg_846 <= _GEN_1870;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_847 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h34f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_847 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_847 <= _GEN_1871;
      end
    end else begin
      lvtReg_847 <= _GEN_1871;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_848 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h350 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_848 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_848 <= _GEN_1872;
      end
    end else begin
      lvtReg_848 <= _GEN_1872;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_849 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h351 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_849 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_849 <= _GEN_1873;
      end
    end else begin
      lvtReg_849 <= _GEN_1873;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_850 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h352 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_850 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_850 <= _GEN_1874;
      end
    end else begin
      lvtReg_850 <= _GEN_1874;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_851 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h353 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_851 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_851 <= _GEN_1875;
      end
    end else begin
      lvtReg_851 <= _GEN_1875;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_852 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h354 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_852 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_852 <= _GEN_1876;
      end
    end else begin
      lvtReg_852 <= _GEN_1876;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_853 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h355 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_853 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_853 <= _GEN_1877;
      end
    end else begin
      lvtReg_853 <= _GEN_1877;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_854 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h356 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_854 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_854 <= _GEN_1878;
      end
    end else begin
      lvtReg_854 <= _GEN_1878;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_855 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h357 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_855 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_855 <= _GEN_1879;
      end
    end else begin
      lvtReg_855 <= _GEN_1879;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_856 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h358 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_856 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_856 <= _GEN_1880;
      end
    end else begin
      lvtReg_856 <= _GEN_1880;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_857 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h359 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_857 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_857 <= _GEN_1881;
      end
    end else begin
      lvtReg_857 <= _GEN_1881;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_858 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_858 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_858 <= _GEN_1882;
      end
    end else begin
      lvtReg_858 <= _GEN_1882;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_859 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_859 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_859 <= _GEN_1883;
      end
    end else begin
      lvtReg_859 <= _GEN_1883;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_860 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_860 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_860 <= _GEN_1884;
      end
    end else begin
      lvtReg_860 <= _GEN_1884;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_861 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_861 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_861 <= _GEN_1885;
      end
    end else begin
      lvtReg_861 <= _GEN_1885;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_862 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_862 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_862 <= _GEN_1886;
      end
    end else begin
      lvtReg_862 <= _GEN_1886;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_863 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h35f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_863 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_863 <= _GEN_1887;
      end
    end else begin
      lvtReg_863 <= _GEN_1887;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_864 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h360 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_864 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_864 <= _GEN_1888;
      end
    end else begin
      lvtReg_864 <= _GEN_1888;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_865 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h361 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_865 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_865 <= _GEN_1889;
      end
    end else begin
      lvtReg_865 <= _GEN_1889;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_866 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h362 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_866 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_866 <= _GEN_1890;
      end
    end else begin
      lvtReg_866 <= _GEN_1890;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_867 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h363 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_867 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_867 <= _GEN_1891;
      end
    end else begin
      lvtReg_867 <= _GEN_1891;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_868 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h364 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_868 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_868 <= _GEN_1892;
      end
    end else begin
      lvtReg_868 <= _GEN_1892;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_869 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h365 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_869 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_869 <= _GEN_1893;
      end
    end else begin
      lvtReg_869 <= _GEN_1893;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_870 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h366 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_870 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_870 <= _GEN_1894;
      end
    end else begin
      lvtReg_870 <= _GEN_1894;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_871 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h367 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_871 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_871 <= _GEN_1895;
      end
    end else begin
      lvtReg_871 <= _GEN_1895;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_872 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h368 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_872 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_872 <= _GEN_1896;
      end
    end else begin
      lvtReg_872 <= _GEN_1896;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_873 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h369 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_873 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_873 <= _GEN_1897;
      end
    end else begin
      lvtReg_873 <= _GEN_1897;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_874 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_874 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_874 <= _GEN_1898;
      end
    end else begin
      lvtReg_874 <= _GEN_1898;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_875 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_875 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_875 <= _GEN_1899;
      end
    end else begin
      lvtReg_875 <= _GEN_1899;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_876 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_876 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_876 <= _GEN_1900;
      end
    end else begin
      lvtReg_876 <= _GEN_1900;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_877 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_877 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_877 <= _GEN_1901;
      end
    end else begin
      lvtReg_877 <= _GEN_1901;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_878 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_878 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_878 <= _GEN_1902;
      end
    end else begin
      lvtReg_878 <= _GEN_1902;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_879 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h36f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_879 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_879 <= _GEN_1903;
      end
    end else begin
      lvtReg_879 <= _GEN_1903;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_880 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h370 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_880 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_880 <= _GEN_1904;
      end
    end else begin
      lvtReg_880 <= _GEN_1904;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_881 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h371 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_881 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_881 <= _GEN_1905;
      end
    end else begin
      lvtReg_881 <= _GEN_1905;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_882 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h372 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_882 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_882 <= _GEN_1906;
      end
    end else begin
      lvtReg_882 <= _GEN_1906;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_883 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h373 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_883 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_883 <= _GEN_1907;
      end
    end else begin
      lvtReg_883 <= _GEN_1907;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_884 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h374 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_884 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_884 <= _GEN_1908;
      end
    end else begin
      lvtReg_884 <= _GEN_1908;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_885 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h375 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_885 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_885 <= _GEN_1909;
      end
    end else begin
      lvtReg_885 <= _GEN_1909;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_886 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h376 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_886 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_886 <= _GEN_1910;
      end
    end else begin
      lvtReg_886 <= _GEN_1910;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_887 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h377 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_887 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_887 <= _GEN_1911;
      end
    end else begin
      lvtReg_887 <= _GEN_1911;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_888 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h378 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_888 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_888 <= _GEN_1912;
      end
    end else begin
      lvtReg_888 <= _GEN_1912;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_889 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h379 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_889 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_889 <= _GEN_1913;
      end
    end else begin
      lvtReg_889 <= _GEN_1913;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_890 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_890 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_890 <= _GEN_1914;
      end
    end else begin
      lvtReg_890 <= _GEN_1914;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_891 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_891 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_891 <= _GEN_1915;
      end
    end else begin
      lvtReg_891 <= _GEN_1915;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_892 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_892 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_892 <= _GEN_1916;
      end
    end else begin
      lvtReg_892 <= _GEN_1916;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_893 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_893 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_893 <= _GEN_1917;
      end
    end else begin
      lvtReg_893 <= _GEN_1917;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_894 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_894 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_894 <= _GEN_1918;
      end
    end else begin
      lvtReg_894 <= _GEN_1918;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_895 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h37f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_895 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_895 <= _GEN_1919;
      end
    end else begin
      lvtReg_895 <= _GEN_1919;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_896 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h380 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_896 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_896 <= _GEN_1920;
      end
    end else begin
      lvtReg_896 <= _GEN_1920;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_897 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h381 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_897 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_897 <= _GEN_1921;
      end
    end else begin
      lvtReg_897 <= _GEN_1921;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_898 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h382 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_898 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_898 <= _GEN_1922;
      end
    end else begin
      lvtReg_898 <= _GEN_1922;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_899 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h383 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_899 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_899 <= _GEN_1923;
      end
    end else begin
      lvtReg_899 <= _GEN_1923;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_900 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h384 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_900 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_900 <= _GEN_1924;
      end
    end else begin
      lvtReg_900 <= _GEN_1924;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_901 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h385 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_901 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_901 <= _GEN_1925;
      end
    end else begin
      lvtReg_901 <= _GEN_1925;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_902 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h386 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_902 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_902 <= _GEN_1926;
      end
    end else begin
      lvtReg_902 <= _GEN_1926;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_903 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h387 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_903 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_903 <= _GEN_1927;
      end
    end else begin
      lvtReg_903 <= _GEN_1927;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_904 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h388 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_904 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_904 <= _GEN_1928;
      end
    end else begin
      lvtReg_904 <= _GEN_1928;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_905 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h389 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_905 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_905 <= _GEN_1929;
      end
    end else begin
      lvtReg_905 <= _GEN_1929;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_906 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_906 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_906 <= _GEN_1930;
      end
    end else begin
      lvtReg_906 <= _GEN_1930;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_907 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_907 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_907 <= _GEN_1931;
      end
    end else begin
      lvtReg_907 <= _GEN_1931;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_908 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_908 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_908 <= _GEN_1932;
      end
    end else begin
      lvtReg_908 <= _GEN_1932;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_909 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_909 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_909 <= _GEN_1933;
      end
    end else begin
      lvtReg_909 <= _GEN_1933;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_910 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_910 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_910 <= _GEN_1934;
      end
    end else begin
      lvtReg_910 <= _GEN_1934;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_911 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h38f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_911 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_911 <= _GEN_1935;
      end
    end else begin
      lvtReg_911 <= _GEN_1935;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_912 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h390 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_912 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_912 <= _GEN_1936;
      end
    end else begin
      lvtReg_912 <= _GEN_1936;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_913 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h391 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_913 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_913 <= _GEN_1937;
      end
    end else begin
      lvtReg_913 <= _GEN_1937;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_914 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h392 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_914 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_914 <= _GEN_1938;
      end
    end else begin
      lvtReg_914 <= _GEN_1938;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_915 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h393 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_915 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_915 <= _GEN_1939;
      end
    end else begin
      lvtReg_915 <= _GEN_1939;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_916 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h394 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_916 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_916 <= _GEN_1940;
      end
    end else begin
      lvtReg_916 <= _GEN_1940;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_917 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h395 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_917 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_917 <= _GEN_1941;
      end
    end else begin
      lvtReg_917 <= _GEN_1941;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_918 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h396 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_918 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_918 <= _GEN_1942;
      end
    end else begin
      lvtReg_918 <= _GEN_1942;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_919 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h397 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_919 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_919 <= _GEN_1943;
      end
    end else begin
      lvtReg_919 <= _GEN_1943;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_920 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h398 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_920 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_920 <= _GEN_1944;
      end
    end else begin
      lvtReg_920 <= _GEN_1944;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_921 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h399 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_921 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_921 <= _GEN_1945;
      end
    end else begin
      lvtReg_921 <= _GEN_1945;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_922 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39a == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_922 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_922 <= _GEN_1946;
      end
    end else begin
      lvtReg_922 <= _GEN_1946;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_923 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39b == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_923 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_923 <= _GEN_1947;
      end
    end else begin
      lvtReg_923 <= _GEN_1947;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_924 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39c == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_924 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_924 <= _GEN_1948;
      end
    end else begin
      lvtReg_924 <= _GEN_1948;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_925 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39d == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_925 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_925 <= _GEN_1949;
      end
    end else begin
      lvtReg_925 <= _GEN_1949;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_926 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39e == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_926 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_926 <= _GEN_1950;
      end
    end else begin
      lvtReg_926 <= _GEN_1950;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_927 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h39f == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_927 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_927 <= _GEN_1951;
      end
    end else begin
      lvtReg_927 <= _GEN_1951;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_928 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_928 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_928 <= _GEN_1952;
      end
    end else begin
      lvtReg_928 <= _GEN_1952;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_929 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_929 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_929 <= _GEN_1953;
      end
    end else begin
      lvtReg_929 <= _GEN_1953;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_930 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_930 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_930 <= _GEN_1954;
      end
    end else begin
      lvtReg_930 <= _GEN_1954;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_931 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_931 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_931 <= _GEN_1955;
      end
    end else begin
      lvtReg_931 <= _GEN_1955;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_932 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_932 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_932 <= _GEN_1956;
      end
    end else begin
      lvtReg_932 <= _GEN_1956;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_933 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_933 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_933 <= _GEN_1957;
      end
    end else begin
      lvtReg_933 <= _GEN_1957;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_934 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_934 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_934 <= _GEN_1958;
      end
    end else begin
      lvtReg_934 <= _GEN_1958;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_935 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_935 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_935 <= _GEN_1959;
      end
    end else begin
      lvtReg_935 <= _GEN_1959;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_936 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_936 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_936 <= _GEN_1960;
      end
    end else begin
      lvtReg_936 <= _GEN_1960;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_937 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3a9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_937 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_937 <= _GEN_1961;
      end
    end else begin
      lvtReg_937 <= _GEN_1961;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_938 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3aa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_938 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_938 <= _GEN_1962;
      end
    end else begin
      lvtReg_938 <= _GEN_1962;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_939 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ab == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_939 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_939 <= _GEN_1963;
      end
    end else begin
      lvtReg_939 <= _GEN_1963;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_940 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ac == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_940 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_940 <= _GEN_1964;
      end
    end else begin
      lvtReg_940 <= _GEN_1964;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_941 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ad == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_941 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_941 <= _GEN_1965;
      end
    end else begin
      lvtReg_941 <= _GEN_1965;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_942 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ae == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_942 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_942 <= _GEN_1966;
      end
    end else begin
      lvtReg_942 <= _GEN_1966;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_943 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3af == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_943 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_943 <= _GEN_1967;
      end
    end else begin
      lvtReg_943 <= _GEN_1967;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_944 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_944 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_944 <= _GEN_1968;
      end
    end else begin
      lvtReg_944 <= _GEN_1968;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_945 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_945 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_945 <= _GEN_1969;
      end
    end else begin
      lvtReg_945 <= _GEN_1969;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_946 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_946 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_946 <= _GEN_1970;
      end
    end else begin
      lvtReg_946 <= _GEN_1970;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_947 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_947 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_947 <= _GEN_1971;
      end
    end else begin
      lvtReg_947 <= _GEN_1971;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_948 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_948 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_948 <= _GEN_1972;
      end
    end else begin
      lvtReg_948 <= _GEN_1972;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_949 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_949 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_949 <= _GEN_1973;
      end
    end else begin
      lvtReg_949 <= _GEN_1973;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_950 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_950 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_950 <= _GEN_1974;
      end
    end else begin
      lvtReg_950 <= _GEN_1974;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_951 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_951 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_951 <= _GEN_1975;
      end
    end else begin
      lvtReg_951 <= _GEN_1975;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_952 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_952 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_952 <= _GEN_1976;
      end
    end else begin
      lvtReg_952 <= _GEN_1976;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_953 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3b9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_953 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_953 <= _GEN_1977;
      end
    end else begin
      lvtReg_953 <= _GEN_1977;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_954 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ba == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_954 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_954 <= _GEN_1978;
      end
    end else begin
      lvtReg_954 <= _GEN_1978;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_955 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3bb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_955 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_955 <= _GEN_1979;
      end
    end else begin
      lvtReg_955 <= _GEN_1979;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_956 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3bc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_956 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_956 <= _GEN_1980;
      end
    end else begin
      lvtReg_956 <= _GEN_1980;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_957 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3bd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_957 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_957 <= _GEN_1981;
      end
    end else begin
      lvtReg_957 <= _GEN_1981;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_958 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3be == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_958 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_958 <= _GEN_1982;
      end
    end else begin
      lvtReg_958 <= _GEN_1982;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_959 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3bf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_959 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_959 <= _GEN_1983;
      end
    end else begin
      lvtReg_959 <= _GEN_1983;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_960 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_960 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_960 <= _GEN_1984;
      end
    end else begin
      lvtReg_960 <= _GEN_1984;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_961 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_961 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_961 <= _GEN_1985;
      end
    end else begin
      lvtReg_961 <= _GEN_1985;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_962 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_962 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_962 <= _GEN_1986;
      end
    end else begin
      lvtReg_962 <= _GEN_1986;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_963 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_963 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_963 <= _GEN_1987;
      end
    end else begin
      lvtReg_963 <= _GEN_1987;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_964 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_964 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_964 <= _GEN_1988;
      end
    end else begin
      lvtReg_964 <= _GEN_1988;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_965 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_965 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_965 <= _GEN_1989;
      end
    end else begin
      lvtReg_965 <= _GEN_1989;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_966 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_966 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_966 <= _GEN_1990;
      end
    end else begin
      lvtReg_966 <= _GEN_1990;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_967 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_967 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_967 <= _GEN_1991;
      end
    end else begin
      lvtReg_967 <= _GEN_1991;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_968 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_968 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_968 <= _GEN_1992;
      end
    end else begin
      lvtReg_968 <= _GEN_1992;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_969 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3c9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_969 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_969 <= _GEN_1993;
      end
    end else begin
      lvtReg_969 <= _GEN_1993;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_970 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ca == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_970 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_970 <= _GEN_1994;
      end
    end else begin
      lvtReg_970 <= _GEN_1994;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_971 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3cb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_971 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_971 <= _GEN_1995;
      end
    end else begin
      lvtReg_971 <= _GEN_1995;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_972 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3cc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_972 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_972 <= _GEN_1996;
      end
    end else begin
      lvtReg_972 <= _GEN_1996;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_973 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3cd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_973 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_973 <= _GEN_1997;
      end
    end else begin
      lvtReg_973 <= _GEN_1997;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_974 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ce == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_974 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_974 <= _GEN_1998;
      end
    end else begin
      lvtReg_974 <= _GEN_1998;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_975 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3cf == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_975 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_975 <= _GEN_1999;
      end
    end else begin
      lvtReg_975 <= _GEN_1999;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_976 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_976 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_976 <= _GEN_2000;
      end
    end else begin
      lvtReg_976 <= _GEN_2000;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_977 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_977 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_977 <= _GEN_2001;
      end
    end else begin
      lvtReg_977 <= _GEN_2001;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_978 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_978 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_978 <= _GEN_2002;
      end
    end else begin
      lvtReg_978 <= _GEN_2002;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_979 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_979 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_979 <= _GEN_2003;
      end
    end else begin
      lvtReg_979 <= _GEN_2003;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_980 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_980 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_980 <= _GEN_2004;
      end
    end else begin
      lvtReg_980 <= _GEN_2004;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_981 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_981 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_981 <= _GEN_2005;
      end
    end else begin
      lvtReg_981 <= _GEN_2005;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_982 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_982 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_982 <= _GEN_2006;
      end
    end else begin
      lvtReg_982 <= _GEN_2006;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_983 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_983 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_983 <= _GEN_2007;
      end
    end else begin
      lvtReg_983 <= _GEN_2007;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_984 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_984 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_984 <= _GEN_2008;
      end
    end else begin
      lvtReg_984 <= _GEN_2008;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_985 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3d9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_985 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_985 <= _GEN_2009;
      end
    end else begin
      lvtReg_985 <= _GEN_2009;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_986 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3da == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_986 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_986 <= _GEN_2010;
      end
    end else begin
      lvtReg_986 <= _GEN_2010;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_987 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3db == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_987 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_987 <= _GEN_2011;
      end
    end else begin
      lvtReg_987 <= _GEN_2011;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_988 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3dc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_988 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_988 <= _GEN_2012;
      end
    end else begin
      lvtReg_988 <= _GEN_2012;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_989 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3dd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_989 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_989 <= _GEN_2013;
      end
    end else begin
      lvtReg_989 <= _GEN_2013;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_990 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3de == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_990 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_990 <= _GEN_2014;
      end
    end else begin
      lvtReg_990 <= _GEN_2014;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_991 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3df == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_991 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_991 <= _GEN_2015;
      end
    end else begin
      lvtReg_991 <= _GEN_2015;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_992 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_992 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_992 <= _GEN_2016;
      end
    end else begin
      lvtReg_992 <= _GEN_2016;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_993 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_993 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_993 <= _GEN_2017;
      end
    end else begin
      lvtReg_993 <= _GEN_2017;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_994 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_994 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_994 <= _GEN_2018;
      end
    end else begin
      lvtReg_994 <= _GEN_2018;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_995 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_995 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_995 <= _GEN_2019;
      end
    end else begin
      lvtReg_995 <= _GEN_2019;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_996 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_996 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_996 <= _GEN_2020;
      end
    end else begin
      lvtReg_996 <= _GEN_2020;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_997 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_997 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_997 <= _GEN_2021;
      end
    end else begin
      lvtReg_997 <= _GEN_2021;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_998 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_998 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_998 <= _GEN_2022;
      end
    end else begin
      lvtReg_998 <= _GEN_2022;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_999 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_999 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_999 <= _GEN_2023;
      end
    end else begin
      lvtReg_999 <= _GEN_2023;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1000 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1000 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1000 <= _GEN_2024;
      end
    end else begin
      lvtReg_1000 <= _GEN_2024;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1001 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3e9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1001 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1001 <= _GEN_2025;
      end
    end else begin
      lvtReg_1001 <= _GEN_2025;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1002 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ea == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1002 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1002 <= _GEN_2026;
      end
    end else begin
      lvtReg_1002 <= _GEN_2026;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1003 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3eb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1003 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1003 <= _GEN_2027;
      end
    end else begin
      lvtReg_1003 <= _GEN_2027;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1004 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ec == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1004 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1004 <= _GEN_2028;
      end
    end else begin
      lvtReg_1004 <= _GEN_2028;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1005 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ed == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1005 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1005 <= _GEN_2029;
      end
    end else begin
      lvtReg_1005 <= _GEN_2029;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1006 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ee == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1006 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1006 <= _GEN_2030;
      end
    end else begin
      lvtReg_1006 <= _GEN_2030;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1007 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ef == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1007 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1007 <= _GEN_2031;
      end
    end else begin
      lvtReg_1007 <= _GEN_2031;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1008 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f0 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1008 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1008 <= _GEN_2032;
      end
    end else begin
      lvtReg_1008 <= _GEN_2032;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1009 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f1 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1009 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1009 <= _GEN_2033;
      end
    end else begin
      lvtReg_1009 <= _GEN_2033;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1010 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f2 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1010 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1010 <= _GEN_2034;
      end
    end else begin
      lvtReg_1010 <= _GEN_2034;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1011 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f3 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1011 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1011 <= _GEN_2035;
      end
    end else begin
      lvtReg_1011 <= _GEN_2035;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1012 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f4 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1012 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1012 <= _GEN_2036;
      end
    end else begin
      lvtReg_1012 <= _GEN_2036;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1013 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f5 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1013 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1013 <= _GEN_2037;
      end
    end else begin
      lvtReg_1013 <= _GEN_2037;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1014 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f6 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1014 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1014 <= _GEN_2038;
      end
    end else begin
      lvtReg_1014 <= _GEN_2038;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1015 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f7 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1015 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1015 <= _GEN_2039;
      end
    end else begin
      lvtReg_1015 <= _GEN_2039;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1016 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f8 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1016 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1016 <= _GEN_2040;
      end
    end else begin
      lvtReg_1016 <= _GEN_2040;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1017 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3f9 == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1017 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1017 <= _GEN_2041;
      end
    end else begin
      lvtReg_1017 <= _GEN_2041;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1018 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3fa == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1018 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1018 <= _GEN_2042;
      end
    end else begin
      lvtReg_1018 <= _GEN_2042;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1019 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3fb == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1019 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1019 <= _GEN_2043;
      end
    end else begin
      lvtReg_1019 <= _GEN_2043;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1020 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3fc == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1020 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1020 <= _GEN_2044;
      end
    end else begin
      lvtReg_1020 <= _GEN_2044;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1021 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3fd == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1021 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1021 <= _GEN_2045;
      end
    end else begin
      lvtReg_1021 <= _GEN_2045;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1022 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3fe == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1022 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1022 <= _GEN_2046;
      end
    end else begin
      lvtReg_1022 <= _GEN_2046;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1023 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (10'h3ff == io_wrAddr_1) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1023 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1023 <= _GEN_2047;
      end
    end else begin
      lvtReg_1023 <= _GEN_2047;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lvtReg_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  lvtReg_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  lvtReg_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  lvtReg_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  lvtReg_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  lvtReg_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  lvtReg_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  lvtReg_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  lvtReg_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  lvtReg_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  lvtReg_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  lvtReg_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  lvtReg_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  lvtReg_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  lvtReg_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  lvtReg_15 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  lvtReg_16 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  lvtReg_17 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  lvtReg_18 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  lvtReg_19 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  lvtReg_20 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  lvtReg_21 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  lvtReg_22 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  lvtReg_23 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  lvtReg_24 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  lvtReg_25 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  lvtReg_26 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  lvtReg_27 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  lvtReg_28 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  lvtReg_29 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  lvtReg_30 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  lvtReg_31 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  lvtReg_32 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  lvtReg_33 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  lvtReg_34 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  lvtReg_35 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  lvtReg_36 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  lvtReg_37 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  lvtReg_38 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  lvtReg_39 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  lvtReg_40 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  lvtReg_41 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  lvtReg_42 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  lvtReg_43 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  lvtReg_44 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  lvtReg_45 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  lvtReg_46 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  lvtReg_47 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  lvtReg_48 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  lvtReg_49 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  lvtReg_50 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  lvtReg_51 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  lvtReg_52 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  lvtReg_53 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  lvtReg_54 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  lvtReg_55 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  lvtReg_56 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  lvtReg_57 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  lvtReg_58 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  lvtReg_59 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  lvtReg_60 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  lvtReg_61 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  lvtReg_62 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  lvtReg_63 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  lvtReg_64 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  lvtReg_65 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  lvtReg_66 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  lvtReg_67 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  lvtReg_68 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  lvtReg_69 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  lvtReg_70 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  lvtReg_71 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  lvtReg_72 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  lvtReg_73 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  lvtReg_74 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  lvtReg_75 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  lvtReg_76 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  lvtReg_77 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  lvtReg_78 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  lvtReg_79 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  lvtReg_80 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  lvtReg_81 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  lvtReg_82 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  lvtReg_83 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  lvtReg_84 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  lvtReg_85 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  lvtReg_86 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  lvtReg_87 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  lvtReg_88 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  lvtReg_89 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  lvtReg_90 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  lvtReg_91 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  lvtReg_92 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  lvtReg_93 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  lvtReg_94 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  lvtReg_95 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  lvtReg_96 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  lvtReg_97 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  lvtReg_98 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  lvtReg_99 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  lvtReg_100 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  lvtReg_101 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  lvtReg_102 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  lvtReg_103 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  lvtReg_104 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  lvtReg_105 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  lvtReg_106 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  lvtReg_107 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  lvtReg_108 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  lvtReg_109 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  lvtReg_110 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  lvtReg_111 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  lvtReg_112 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  lvtReg_113 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  lvtReg_114 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  lvtReg_115 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  lvtReg_116 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  lvtReg_117 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  lvtReg_118 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  lvtReg_119 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  lvtReg_120 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  lvtReg_121 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  lvtReg_122 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  lvtReg_123 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  lvtReg_124 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  lvtReg_125 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  lvtReg_126 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  lvtReg_127 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  lvtReg_128 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  lvtReg_129 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  lvtReg_130 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  lvtReg_131 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  lvtReg_132 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  lvtReg_133 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  lvtReg_134 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  lvtReg_135 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  lvtReg_136 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  lvtReg_137 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  lvtReg_138 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  lvtReg_139 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  lvtReg_140 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  lvtReg_141 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  lvtReg_142 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  lvtReg_143 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  lvtReg_144 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  lvtReg_145 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  lvtReg_146 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  lvtReg_147 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  lvtReg_148 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  lvtReg_149 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  lvtReg_150 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  lvtReg_151 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  lvtReg_152 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  lvtReg_153 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  lvtReg_154 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  lvtReg_155 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  lvtReg_156 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  lvtReg_157 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  lvtReg_158 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  lvtReg_159 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  lvtReg_160 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  lvtReg_161 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  lvtReg_162 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  lvtReg_163 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  lvtReg_164 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  lvtReg_165 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  lvtReg_166 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  lvtReg_167 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  lvtReg_168 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  lvtReg_169 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  lvtReg_170 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  lvtReg_171 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  lvtReg_172 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  lvtReg_173 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  lvtReg_174 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  lvtReg_175 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  lvtReg_176 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  lvtReg_177 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  lvtReg_178 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  lvtReg_179 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  lvtReg_180 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  lvtReg_181 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  lvtReg_182 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  lvtReg_183 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  lvtReg_184 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  lvtReg_185 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  lvtReg_186 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  lvtReg_187 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  lvtReg_188 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  lvtReg_189 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  lvtReg_190 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  lvtReg_191 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  lvtReg_192 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  lvtReg_193 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  lvtReg_194 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  lvtReg_195 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  lvtReg_196 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  lvtReg_197 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  lvtReg_198 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  lvtReg_199 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  lvtReg_200 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  lvtReg_201 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  lvtReg_202 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  lvtReg_203 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  lvtReg_204 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  lvtReg_205 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  lvtReg_206 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  lvtReg_207 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  lvtReg_208 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  lvtReg_209 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  lvtReg_210 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  lvtReg_211 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  lvtReg_212 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  lvtReg_213 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  lvtReg_214 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  lvtReg_215 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  lvtReg_216 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  lvtReg_217 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  lvtReg_218 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  lvtReg_219 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  lvtReg_220 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  lvtReg_221 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  lvtReg_222 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  lvtReg_223 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  lvtReg_224 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  lvtReg_225 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  lvtReg_226 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  lvtReg_227 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  lvtReg_228 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  lvtReg_229 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  lvtReg_230 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  lvtReg_231 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  lvtReg_232 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  lvtReg_233 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  lvtReg_234 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  lvtReg_235 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  lvtReg_236 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  lvtReg_237 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  lvtReg_238 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  lvtReg_239 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  lvtReg_240 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  lvtReg_241 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  lvtReg_242 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  lvtReg_243 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  lvtReg_244 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  lvtReg_245 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  lvtReg_246 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  lvtReg_247 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  lvtReg_248 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  lvtReg_249 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  lvtReg_250 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  lvtReg_251 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  lvtReg_252 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  lvtReg_253 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  lvtReg_254 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  lvtReg_255 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  lvtReg_256 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  lvtReg_257 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  lvtReg_258 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  lvtReg_259 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  lvtReg_260 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  lvtReg_261 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  lvtReg_262 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  lvtReg_263 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  lvtReg_264 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  lvtReg_265 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  lvtReg_266 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  lvtReg_267 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  lvtReg_268 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  lvtReg_269 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  lvtReg_270 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  lvtReg_271 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  lvtReg_272 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  lvtReg_273 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  lvtReg_274 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  lvtReg_275 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  lvtReg_276 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  lvtReg_277 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  lvtReg_278 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  lvtReg_279 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  lvtReg_280 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  lvtReg_281 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  lvtReg_282 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  lvtReg_283 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  lvtReg_284 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  lvtReg_285 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  lvtReg_286 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  lvtReg_287 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  lvtReg_288 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  lvtReg_289 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  lvtReg_290 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  lvtReg_291 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  lvtReg_292 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  lvtReg_293 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  lvtReg_294 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  lvtReg_295 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  lvtReg_296 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  lvtReg_297 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  lvtReg_298 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  lvtReg_299 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  lvtReg_300 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  lvtReg_301 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  lvtReg_302 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  lvtReg_303 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  lvtReg_304 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  lvtReg_305 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  lvtReg_306 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  lvtReg_307 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  lvtReg_308 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  lvtReg_309 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  lvtReg_310 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  lvtReg_311 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  lvtReg_312 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  lvtReg_313 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  lvtReg_314 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  lvtReg_315 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  lvtReg_316 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  lvtReg_317 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  lvtReg_318 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  lvtReg_319 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  lvtReg_320 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  lvtReg_321 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  lvtReg_322 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  lvtReg_323 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  lvtReg_324 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  lvtReg_325 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  lvtReg_326 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  lvtReg_327 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  lvtReg_328 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  lvtReg_329 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  lvtReg_330 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  lvtReg_331 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  lvtReg_332 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  lvtReg_333 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  lvtReg_334 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  lvtReg_335 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  lvtReg_336 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  lvtReg_337 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  lvtReg_338 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  lvtReg_339 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  lvtReg_340 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  lvtReg_341 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  lvtReg_342 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  lvtReg_343 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  lvtReg_344 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  lvtReg_345 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  lvtReg_346 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  lvtReg_347 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  lvtReg_348 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  lvtReg_349 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  lvtReg_350 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  lvtReg_351 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  lvtReg_352 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  lvtReg_353 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  lvtReg_354 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  lvtReg_355 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  lvtReg_356 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  lvtReg_357 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  lvtReg_358 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  lvtReg_359 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  lvtReg_360 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  lvtReg_361 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  lvtReg_362 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  lvtReg_363 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  lvtReg_364 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  lvtReg_365 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  lvtReg_366 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  lvtReg_367 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  lvtReg_368 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  lvtReg_369 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  lvtReg_370 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  lvtReg_371 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  lvtReg_372 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  lvtReg_373 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  lvtReg_374 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  lvtReg_375 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  lvtReg_376 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  lvtReg_377 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  lvtReg_378 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  lvtReg_379 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  lvtReg_380 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  lvtReg_381 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  lvtReg_382 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  lvtReg_383 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  lvtReg_384 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  lvtReg_385 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  lvtReg_386 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  lvtReg_387 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  lvtReg_388 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  lvtReg_389 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  lvtReg_390 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  lvtReg_391 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  lvtReg_392 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  lvtReg_393 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  lvtReg_394 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  lvtReg_395 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  lvtReg_396 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  lvtReg_397 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  lvtReg_398 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  lvtReg_399 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  lvtReg_400 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  lvtReg_401 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  lvtReg_402 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  lvtReg_403 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  lvtReg_404 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  lvtReg_405 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  lvtReg_406 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  lvtReg_407 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  lvtReg_408 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  lvtReg_409 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  lvtReg_410 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  lvtReg_411 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  lvtReg_412 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  lvtReg_413 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  lvtReg_414 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  lvtReg_415 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  lvtReg_416 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  lvtReg_417 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  lvtReg_418 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  lvtReg_419 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  lvtReg_420 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  lvtReg_421 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  lvtReg_422 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  lvtReg_423 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  lvtReg_424 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  lvtReg_425 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  lvtReg_426 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  lvtReg_427 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  lvtReg_428 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  lvtReg_429 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  lvtReg_430 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  lvtReg_431 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  lvtReg_432 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  lvtReg_433 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  lvtReg_434 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  lvtReg_435 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  lvtReg_436 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  lvtReg_437 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  lvtReg_438 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  lvtReg_439 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  lvtReg_440 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  lvtReg_441 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  lvtReg_442 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  lvtReg_443 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  lvtReg_444 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  lvtReg_445 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  lvtReg_446 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  lvtReg_447 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  lvtReg_448 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  lvtReg_449 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  lvtReg_450 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  lvtReg_451 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  lvtReg_452 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  lvtReg_453 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  lvtReg_454 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  lvtReg_455 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  lvtReg_456 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  lvtReg_457 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  lvtReg_458 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  lvtReg_459 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  lvtReg_460 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  lvtReg_461 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  lvtReg_462 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  lvtReg_463 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  lvtReg_464 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  lvtReg_465 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  lvtReg_466 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  lvtReg_467 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  lvtReg_468 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  lvtReg_469 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  lvtReg_470 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  lvtReg_471 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  lvtReg_472 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  lvtReg_473 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  lvtReg_474 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  lvtReg_475 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  lvtReg_476 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  lvtReg_477 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  lvtReg_478 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  lvtReg_479 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  lvtReg_480 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  lvtReg_481 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  lvtReg_482 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  lvtReg_483 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  lvtReg_484 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  lvtReg_485 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  lvtReg_486 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  lvtReg_487 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  lvtReg_488 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  lvtReg_489 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  lvtReg_490 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  lvtReg_491 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  lvtReg_492 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  lvtReg_493 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  lvtReg_494 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  lvtReg_495 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  lvtReg_496 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  lvtReg_497 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  lvtReg_498 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  lvtReg_499 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  lvtReg_500 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  lvtReg_501 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  lvtReg_502 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  lvtReg_503 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  lvtReg_504 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  lvtReg_505 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  lvtReg_506 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  lvtReg_507 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  lvtReg_508 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  lvtReg_509 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  lvtReg_510 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  lvtReg_511 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  lvtReg_512 = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  lvtReg_513 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  lvtReg_514 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  lvtReg_515 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  lvtReg_516 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  lvtReg_517 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  lvtReg_518 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  lvtReg_519 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  lvtReg_520 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  lvtReg_521 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  lvtReg_522 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  lvtReg_523 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  lvtReg_524 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  lvtReg_525 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  lvtReg_526 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  lvtReg_527 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  lvtReg_528 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  lvtReg_529 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  lvtReg_530 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  lvtReg_531 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  lvtReg_532 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  lvtReg_533 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  lvtReg_534 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  lvtReg_535 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  lvtReg_536 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  lvtReg_537 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  lvtReg_538 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  lvtReg_539 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  lvtReg_540 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  lvtReg_541 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  lvtReg_542 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  lvtReg_543 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  lvtReg_544 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  lvtReg_545 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  lvtReg_546 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  lvtReg_547 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  lvtReg_548 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  lvtReg_549 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  lvtReg_550 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  lvtReg_551 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  lvtReg_552 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  lvtReg_553 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  lvtReg_554 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  lvtReg_555 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  lvtReg_556 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  lvtReg_557 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  lvtReg_558 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  lvtReg_559 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  lvtReg_560 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  lvtReg_561 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  lvtReg_562 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  lvtReg_563 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  lvtReg_564 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  lvtReg_565 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  lvtReg_566 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  lvtReg_567 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  lvtReg_568 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  lvtReg_569 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  lvtReg_570 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  lvtReg_571 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  lvtReg_572 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  lvtReg_573 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  lvtReg_574 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  lvtReg_575 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  lvtReg_576 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  lvtReg_577 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  lvtReg_578 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  lvtReg_579 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  lvtReg_580 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  lvtReg_581 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  lvtReg_582 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  lvtReg_583 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  lvtReg_584 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  lvtReg_585 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  lvtReg_586 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  lvtReg_587 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  lvtReg_588 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  lvtReg_589 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  lvtReg_590 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  lvtReg_591 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  lvtReg_592 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  lvtReg_593 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  lvtReg_594 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  lvtReg_595 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  lvtReg_596 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  lvtReg_597 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  lvtReg_598 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  lvtReg_599 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  lvtReg_600 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  lvtReg_601 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  lvtReg_602 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  lvtReg_603 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  lvtReg_604 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  lvtReg_605 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  lvtReg_606 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  lvtReg_607 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  lvtReg_608 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  lvtReg_609 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  lvtReg_610 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  lvtReg_611 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  lvtReg_612 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  lvtReg_613 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  lvtReg_614 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  lvtReg_615 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  lvtReg_616 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  lvtReg_617 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  lvtReg_618 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  lvtReg_619 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  lvtReg_620 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  lvtReg_621 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  lvtReg_622 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  lvtReg_623 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  lvtReg_624 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  lvtReg_625 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  lvtReg_626 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  lvtReg_627 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  lvtReg_628 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  lvtReg_629 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  lvtReg_630 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  lvtReg_631 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  lvtReg_632 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  lvtReg_633 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  lvtReg_634 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  lvtReg_635 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  lvtReg_636 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  lvtReg_637 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  lvtReg_638 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  lvtReg_639 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  lvtReg_640 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  lvtReg_641 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  lvtReg_642 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  lvtReg_643 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  lvtReg_644 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  lvtReg_645 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  lvtReg_646 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  lvtReg_647 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  lvtReg_648 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  lvtReg_649 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  lvtReg_650 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  lvtReg_651 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  lvtReg_652 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  lvtReg_653 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  lvtReg_654 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  lvtReg_655 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  lvtReg_656 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  lvtReg_657 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  lvtReg_658 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  lvtReg_659 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  lvtReg_660 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  lvtReg_661 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  lvtReg_662 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  lvtReg_663 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  lvtReg_664 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  lvtReg_665 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  lvtReg_666 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  lvtReg_667 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  lvtReg_668 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  lvtReg_669 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  lvtReg_670 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  lvtReg_671 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  lvtReg_672 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  lvtReg_673 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  lvtReg_674 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  lvtReg_675 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  lvtReg_676 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  lvtReg_677 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  lvtReg_678 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  lvtReg_679 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  lvtReg_680 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  lvtReg_681 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  lvtReg_682 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  lvtReg_683 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  lvtReg_684 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  lvtReg_685 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  lvtReg_686 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  lvtReg_687 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  lvtReg_688 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  lvtReg_689 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  lvtReg_690 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  lvtReg_691 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  lvtReg_692 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  lvtReg_693 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  lvtReg_694 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  lvtReg_695 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  lvtReg_696 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  lvtReg_697 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  lvtReg_698 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  lvtReg_699 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  lvtReg_700 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  lvtReg_701 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  lvtReg_702 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  lvtReg_703 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  lvtReg_704 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  lvtReg_705 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  lvtReg_706 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  lvtReg_707 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  lvtReg_708 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  lvtReg_709 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  lvtReg_710 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  lvtReg_711 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  lvtReg_712 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  lvtReg_713 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  lvtReg_714 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  lvtReg_715 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  lvtReg_716 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  lvtReg_717 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  lvtReg_718 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  lvtReg_719 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  lvtReg_720 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  lvtReg_721 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  lvtReg_722 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  lvtReg_723 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  lvtReg_724 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  lvtReg_725 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  lvtReg_726 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  lvtReg_727 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  lvtReg_728 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  lvtReg_729 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  lvtReg_730 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  lvtReg_731 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  lvtReg_732 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  lvtReg_733 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  lvtReg_734 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  lvtReg_735 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  lvtReg_736 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  lvtReg_737 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  lvtReg_738 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  lvtReg_739 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  lvtReg_740 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  lvtReg_741 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  lvtReg_742 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  lvtReg_743 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  lvtReg_744 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  lvtReg_745 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  lvtReg_746 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  lvtReg_747 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  lvtReg_748 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  lvtReg_749 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  lvtReg_750 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  lvtReg_751 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  lvtReg_752 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  lvtReg_753 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  lvtReg_754 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  lvtReg_755 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  lvtReg_756 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  lvtReg_757 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  lvtReg_758 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  lvtReg_759 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  lvtReg_760 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  lvtReg_761 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  lvtReg_762 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  lvtReg_763 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  lvtReg_764 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  lvtReg_765 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  lvtReg_766 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  lvtReg_767 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  lvtReg_768 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  lvtReg_769 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  lvtReg_770 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  lvtReg_771 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  lvtReg_772 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  lvtReg_773 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  lvtReg_774 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  lvtReg_775 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  lvtReg_776 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  lvtReg_777 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  lvtReg_778 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  lvtReg_779 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  lvtReg_780 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  lvtReg_781 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  lvtReg_782 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  lvtReg_783 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  lvtReg_784 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  lvtReg_785 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  lvtReg_786 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  lvtReg_787 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  lvtReg_788 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  lvtReg_789 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  lvtReg_790 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  lvtReg_791 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  lvtReg_792 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  lvtReg_793 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  lvtReg_794 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  lvtReg_795 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  lvtReg_796 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  lvtReg_797 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  lvtReg_798 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  lvtReg_799 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  lvtReg_800 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  lvtReg_801 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  lvtReg_802 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  lvtReg_803 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  lvtReg_804 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  lvtReg_805 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  lvtReg_806 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  lvtReg_807 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  lvtReg_808 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  lvtReg_809 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  lvtReg_810 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  lvtReg_811 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  lvtReg_812 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  lvtReg_813 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  lvtReg_814 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  lvtReg_815 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  lvtReg_816 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  lvtReg_817 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  lvtReg_818 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  lvtReg_819 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  lvtReg_820 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  lvtReg_821 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  lvtReg_822 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  lvtReg_823 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  lvtReg_824 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  lvtReg_825 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  lvtReg_826 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  lvtReg_827 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  lvtReg_828 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  lvtReg_829 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  lvtReg_830 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  lvtReg_831 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  lvtReg_832 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  lvtReg_833 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  lvtReg_834 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  lvtReg_835 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  lvtReg_836 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  lvtReg_837 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  lvtReg_838 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  lvtReg_839 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  lvtReg_840 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  lvtReg_841 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  lvtReg_842 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  lvtReg_843 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  lvtReg_844 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  lvtReg_845 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  lvtReg_846 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  lvtReg_847 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  lvtReg_848 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  lvtReg_849 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  lvtReg_850 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  lvtReg_851 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  lvtReg_852 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  lvtReg_853 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  lvtReg_854 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  lvtReg_855 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  lvtReg_856 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  lvtReg_857 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  lvtReg_858 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  lvtReg_859 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  lvtReg_860 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  lvtReg_861 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  lvtReg_862 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  lvtReg_863 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  lvtReg_864 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  lvtReg_865 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  lvtReg_866 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  lvtReg_867 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  lvtReg_868 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  lvtReg_869 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  lvtReg_870 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  lvtReg_871 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  lvtReg_872 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  lvtReg_873 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  lvtReg_874 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  lvtReg_875 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  lvtReg_876 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  lvtReg_877 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  lvtReg_878 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  lvtReg_879 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  lvtReg_880 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  lvtReg_881 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  lvtReg_882 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  lvtReg_883 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  lvtReg_884 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  lvtReg_885 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  lvtReg_886 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  lvtReg_887 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  lvtReg_888 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  lvtReg_889 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  lvtReg_890 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  lvtReg_891 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  lvtReg_892 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  lvtReg_893 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  lvtReg_894 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  lvtReg_895 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  lvtReg_896 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  lvtReg_897 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  lvtReg_898 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  lvtReg_899 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  lvtReg_900 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  lvtReg_901 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  lvtReg_902 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  lvtReg_903 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  lvtReg_904 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  lvtReg_905 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  lvtReg_906 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  lvtReg_907 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  lvtReg_908 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  lvtReg_909 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  lvtReg_910 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  lvtReg_911 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  lvtReg_912 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  lvtReg_913 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  lvtReg_914 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  lvtReg_915 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  lvtReg_916 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  lvtReg_917 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  lvtReg_918 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  lvtReg_919 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  lvtReg_920 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  lvtReg_921 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  lvtReg_922 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  lvtReg_923 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  lvtReg_924 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  lvtReg_925 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  lvtReg_926 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  lvtReg_927 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  lvtReg_928 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  lvtReg_929 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  lvtReg_930 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  lvtReg_931 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  lvtReg_932 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  lvtReg_933 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  lvtReg_934 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  lvtReg_935 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  lvtReg_936 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  lvtReg_937 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  lvtReg_938 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  lvtReg_939 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  lvtReg_940 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  lvtReg_941 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  lvtReg_942 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  lvtReg_943 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  lvtReg_944 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  lvtReg_945 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  lvtReg_946 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  lvtReg_947 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  lvtReg_948 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  lvtReg_949 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  lvtReg_950 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  lvtReg_951 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  lvtReg_952 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  lvtReg_953 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  lvtReg_954 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  lvtReg_955 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  lvtReg_956 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  lvtReg_957 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  lvtReg_958 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  lvtReg_959 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  lvtReg_960 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  lvtReg_961 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  lvtReg_962 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  lvtReg_963 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  lvtReg_964 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  lvtReg_965 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  lvtReg_966 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  lvtReg_967 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  lvtReg_968 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  lvtReg_969 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  lvtReg_970 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  lvtReg_971 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  lvtReg_972 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  lvtReg_973 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  lvtReg_974 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  lvtReg_975 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  lvtReg_976 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  lvtReg_977 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  lvtReg_978 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  lvtReg_979 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  lvtReg_980 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  lvtReg_981 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  lvtReg_982 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  lvtReg_983 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  lvtReg_984 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  lvtReg_985 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  lvtReg_986 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  lvtReg_987 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  lvtReg_988 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  lvtReg_989 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  lvtReg_990 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  lvtReg_991 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  lvtReg_992 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  lvtReg_993 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  lvtReg_994 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  lvtReg_995 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  lvtReg_996 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  lvtReg_997 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  lvtReg_998 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  lvtReg_999 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  lvtReg_1000 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  lvtReg_1001 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  lvtReg_1002 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  lvtReg_1003 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  lvtReg_1004 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  lvtReg_1005 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  lvtReg_1006 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  lvtReg_1007 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  lvtReg_1008 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  lvtReg_1009 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  lvtReg_1010 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  lvtReg_1011 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  lvtReg_1012 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  lvtReg_1013 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  lvtReg_1014 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  lvtReg_1015 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  lvtReg_1016 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  lvtReg_1017 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  lvtReg_1018 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  lvtReg_1019 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  lvtReg_1020 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  lvtReg_1021 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  lvtReg_1022 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  lvtReg_1023 = _RAND_1023[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LVTMultiPortRams(
  input        clock,
  input        reset,
  input  [9:0] io_wrAddr_0,
  input  [9:0] io_wrAddr_1,
  input  [7:0] io_wrData_0,
  input  [7:0] io_wrData_1,
  input        io_wrEna_0,
  input        io_wrEna_1,
  input  [9:0] io_rdAddr_0,
  input  [9:0] io_rdAddr_1,
  output [7:0] io_rdData_0,
  output [7:0] io_rdData_1
);
  wire  Memory_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_1_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_1_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_1_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_1_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_1_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_1_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_2_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_2_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_2_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_2_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_2_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_2_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_3_clock; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_3_io_rdAddr; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_3_io_rdData; // @[LVTMultiPortRams.scala 52:44]
  wire  Memory_3_io_wrEna; // @[LVTMultiPortRams.scala 52:44]
  wire [7:0] Memory_3_io_wrData; // @[LVTMultiPortRams.scala 52:44]
  wire [9:0] Memory_3_io_wrAddr; // @[LVTMultiPortRams.scala 52:44]
  wire  lvt_clock; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_reset; // @[LVTMultiPortRams.scala 53:19]
  wire [9:0] lvt_io_wrAddr_0; // @[LVTMultiPortRams.scala 53:19]
  wire [9:0] lvt_io_wrAddr_1; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_io_wrEna_0; // @[LVTMultiPortRams.scala 53:19]
  wire  lvt_io_wrEna_1; // @[LVTMultiPortRams.scala 53:19]
  wire [9:0] lvt_io_rdAddr_0; // @[LVTMultiPortRams.scala 53:19]
  wire [9:0] lvt_io_rdAddr_1; // @[LVTMultiPortRams.scala 53:19]
  wire [1:0] lvt_io_rdIdx_0; // @[LVTMultiPortRams.scala 53:19]
  wire [1:0] lvt_io_rdIdx_1; // @[LVTMultiPortRams.scala 53:19]
  wire [3:0] _io_rdData_0_T = lvt_io_rdIdx_0 * 2'h2; // @[LVTMultiPortRams.scala 72:30]
  wire [4:0] _io_rdData_0_T_1 = {{1'd0}, _io_rdData_0_T}; // @[LVTMultiPortRams.scala 72:36]
  wire [7:0] mems_0_rdData = Memory_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] mems_1_rdData = Memory_1_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_6 = 2'h1 == _io_rdData_0_T_1[1:0] ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_2_rdData = Memory_2_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [7:0] _GEN_11 = 2'h2 == _io_rdData_0_T_1[1:0] ? mems_2_rdData : _GEN_6; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] mems_3_rdData = Memory_3_io_rdData; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 52:21]
  wire [3:0] _io_rdData_1_T = lvt_io_rdIdx_1 * 2'h2; // @[LVTMultiPortRams.scala 72:30]
  wire [3:0] _io_rdData_1_T_2 = _io_rdData_1_T + 4'h1; // @[LVTMultiPortRams.scala 72:36]
  wire [7:0] _GEN_26 = 2'h1 == _io_rdData_1_T_2[1:0] ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  wire [7:0] _GEN_31 = 2'h2 == _io_rdData_1_T_2[1:0] ? mems_2_rdData : _GEN_26; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  Memory Memory ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_clock),
    .io_rdAddr(Memory_io_rdAddr),
    .io_rdData(Memory_io_rdData),
    .io_wrEna(Memory_io_wrEna),
    .io_wrData(Memory_io_wrData),
    .io_wrAddr(Memory_io_wrAddr)
  );
  Memory Memory_1 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_1_clock),
    .io_rdAddr(Memory_1_io_rdAddr),
    .io_rdData(Memory_1_io_rdData),
    .io_wrEna(Memory_1_io_wrEna),
    .io_wrData(Memory_1_io_wrData),
    .io_wrAddr(Memory_1_io_wrAddr)
  );
  Memory Memory_2 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_2_clock),
    .io_rdAddr(Memory_2_io_rdAddr),
    .io_rdData(Memory_2_io_rdData),
    .io_wrEna(Memory_2_io_wrEna),
    .io_wrData(Memory_2_io_wrData),
    .io_wrAddr(Memory_2_io_wrAddr)
  );
  Memory Memory_3 ( // @[LVTMultiPortRams.scala 52:44]
    .clock(Memory_3_clock),
    .io_rdAddr(Memory_3_io_rdAddr),
    .io_rdData(Memory_3_io_rdData),
    .io_wrEna(Memory_3_io_wrEna),
    .io_wrData(Memory_3_io_wrData),
    .io_wrAddr(Memory_3_io_wrAddr)
  );
  LiveValueTable lvt ( // @[LVTMultiPortRams.scala 53:19]
    .clock(lvt_clock),
    .reset(lvt_reset),
    .io_wrAddr_0(lvt_io_wrAddr_0),
    .io_wrAddr_1(lvt_io_wrAddr_1),
    .io_wrEna_0(lvt_io_wrEna_0),
    .io_wrEna_1(lvt_io_wrEna_1),
    .io_rdAddr_0(lvt_io_rdAddr_0),
    .io_rdAddr_1(lvt_io_rdAddr_1),
    .io_rdIdx_0(lvt_io_rdIdx_0),
    .io_rdIdx_1(lvt_io_rdIdx_1)
  );
  assign io_rdData_0 = 2'h3 == _io_rdData_0_T_1[1:0] ? mems_3_rdData : _GEN_11; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  assign io_rdData_1 = 2'h3 == _io_rdData_1_T_2[1:0] ? mems_3_rdData : _GEN_31; // @[LVTMultiPortRams.scala 72:18 LVTMultiPortRams.scala 72:18]
  assign Memory_clock = clock;
  assign Memory_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_1_clock = clock;
  assign Memory_1_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_1_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_1_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_1_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_2_clock = clock;
  assign Memory_2_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_2_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_2_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_2_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign Memory_3_clock = clock;
  assign Memory_3_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 60:30]
  assign Memory_3_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 57:29]
  assign Memory_3_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 59:30]
  assign Memory_3_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 52:21 LVTMultiPortRams.scala 58:30]
  assign lvt_clock = clock;
  assign lvt_reset = reset;
  assign lvt_io_wrAddr_0 = io_wrAddr_0; // @[LVTMultiPortRams.scala 65:22]
  assign lvt_io_wrAddr_1 = io_wrAddr_1; // @[LVTMultiPortRams.scala 65:22]
  assign lvt_io_wrEna_0 = io_wrEna_0; // @[LVTMultiPortRams.scala 64:21]
  assign lvt_io_wrEna_1 = io_wrEna_1; // @[LVTMultiPortRams.scala 64:21]
  assign lvt_io_rdAddr_0 = io_rdAddr_0; // @[LVTMultiPortRams.scala 68:22]
  assign lvt_io_rdAddr_1 = io_rdAddr_1; // @[LVTMultiPortRams.scala 68:22]
endmodule
