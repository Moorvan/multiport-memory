module Memory(
  input        clock,
  input  [9:0] io_rdAddr,
  output [7:0] io_rdData,
  input        io_wrEna,
  input  [7:0] io_wrData,
  input  [9:0] io_wrAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:1023]; // @[Memory.scala 16:24]
  wire [7:0] mem_memData_data; // @[Memory.scala 16:24]
  wire [9:0] mem_memData_addr; // @[Memory.scala 16:24]
  wire [7:0] mem_MPORT_data; // @[Memory.scala 16:24]
  wire [9:0] mem_MPORT_addr; // @[Memory.scala 16:24]
  wire  mem_MPORT_mask; // @[Memory.scala 16:24]
  wire  mem_MPORT_en; // @[Memory.scala 16:24]
  reg [9:0] mem_memData_addr_pipe_0;
  reg [7:0] wrDateReg; // @[Memory.scala 18:26]
  reg  doForwardReg; // @[Memory.scala 19:29]
  assign mem_memData_addr = mem_memData_addr_pipe_0;
  assign mem_memData_data = mem[mem_memData_addr]; // @[Memory.scala 16:24]
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = doForwardReg ? wrDateReg : mem_memData_data; // @[Memory.scala 25:19]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 16:24]
    end
    mem_memData_addr_pipe_0 <= io_rdAddr;
    wrDateReg <= io_wrData; // @[Memory.scala 18:26]
    doForwardReg <= io_wrAddr == io_rdAddr & io_wrEna; // @[Memory.scala 19:54]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_memData_addr_pipe_0 = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  wrDateReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  doForwardReg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LiveValueTable(
  input        clock,
  input        reset,
  input  [9:0] io_wrAddr_0,
  input  [9:0] io_wrAddr_1,
  input        io_wrEna_0,
  input        io_wrEna_1,
  input  [9:0] io_rdAddr_0,
  input  [9:0] io_rdAddr_1,
  output [1:0] io_rdIdx_0,
  output [1:0] io_rdIdx_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] lvtReg_0; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_1; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_2; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_3; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_4; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_5; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_6; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_7; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_8; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_9; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_10; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_11; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_12; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_13; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_14; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_15; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_16; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_17; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_18; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_19; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_20; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_21; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_22; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_23; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_24; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_25; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_26; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_27; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_28; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_29; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_30; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_31; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_32; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_33; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_34; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_35; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_36; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_37; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_38; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_39; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_40; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_41; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_42; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_43; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_44; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_45; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_46; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_47; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_48; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_49; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_50; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_51; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_52; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_53; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_54; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_55; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_56; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_57; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_58; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_59; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_60; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_61; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_62; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_63; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_64; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_65; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_66; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_67; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_68; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_69; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_70; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_71; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_72; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_73; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_74; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_75; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_76; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_77; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_78; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_79; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_80; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_81; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_82; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_83; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_84; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_85; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_86; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_87; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_88; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_89; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_90; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_91; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_92; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_93; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_94; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_95; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_96; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_97; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_98; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_99; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_100; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_101; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_102; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_103; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_104; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_105; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_106; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_107; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_108; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_109; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_110; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_111; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_112; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_113; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_114; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_115; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_116; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_117; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_118; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_119; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_120; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_121; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_122; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_123; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_124; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_125; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_126; // @[LVTMultiPortRams.scala 28:23]
  reg [1:0] lvtReg_127; // @[LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_0 = 7'h0 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_0; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_1 = 7'h1 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_1; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_2 = 7'h2 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_2; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_3 = 7'h3 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_3; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_4 = 7'h4 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_4; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_5 = 7'h5 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_5; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_6 = 7'h6 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_6; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_7 = 7'h7 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_7; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_8 = 7'h8 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_8; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_9 = 7'h9 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_9; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_10 = 7'ha == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_10; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_11 = 7'hb == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_11; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_12 = 7'hc == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_12; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_13 = 7'hd == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_13; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_14 = 7'he == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_14; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_15 = 7'hf == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_15; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_16 = 7'h10 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_16; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_17 = 7'h11 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_17; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_18 = 7'h12 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_18; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_19 = 7'h13 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_19; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_20 = 7'h14 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_20; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_21 = 7'h15 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_21; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_22 = 7'h16 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_22; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_23 = 7'h17 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_23; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_24 = 7'h18 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_24; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_25 = 7'h19 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_25; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_26 = 7'h1a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_26; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_27 = 7'h1b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_27; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_28 = 7'h1c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_28; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_29 = 7'h1d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_29; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_30 = 7'h1e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_30; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_31 = 7'h1f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_31; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_32 = 7'h20 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_32; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_33 = 7'h21 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_33; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_34 = 7'h22 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_34; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_35 = 7'h23 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_35; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_36 = 7'h24 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_36; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_37 = 7'h25 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_37; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_38 = 7'h26 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_38; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_39 = 7'h27 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_39; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_40 = 7'h28 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_40; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_41 = 7'h29 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_41; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_42 = 7'h2a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_42; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_43 = 7'h2b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_43; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_44 = 7'h2c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_44; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_45 = 7'h2d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_45; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_46 = 7'h2e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_46; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_47 = 7'h2f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_47; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_48 = 7'h30 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_48; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_49 = 7'h31 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_49; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_50 = 7'h32 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_50; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_51 = 7'h33 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_51; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_52 = 7'h34 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_52; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_53 = 7'h35 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_53; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_54 = 7'h36 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_54; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_55 = 7'h37 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_55; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_56 = 7'h38 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_56; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_57 = 7'h39 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_57; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_58 = 7'h3a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_58; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_59 = 7'h3b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_59; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_60 = 7'h3c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_60; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_61 = 7'h3d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_61; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_62 = 7'h3e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_62; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_63 = 7'h3f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_63; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_64 = 7'h40 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_64; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_65 = 7'h41 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_65; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_66 = 7'h42 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_66; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_67 = 7'h43 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_67; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_68 = 7'h44 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_68; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_69 = 7'h45 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_69; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_70 = 7'h46 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_70; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_71 = 7'h47 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_71; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_72 = 7'h48 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_72; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_73 = 7'h49 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_73; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_74 = 7'h4a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_74; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_75 = 7'h4b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_75; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_76 = 7'h4c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_76; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_77 = 7'h4d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_77; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_78 = 7'h4e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_78; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_79 = 7'h4f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_79; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_80 = 7'h50 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_80; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_81 = 7'h51 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_81; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_82 = 7'h52 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_82; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_83 = 7'h53 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_83; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_84 = 7'h54 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_84; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_85 = 7'h55 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_85; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_86 = 7'h56 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_86; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_87 = 7'h57 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_87; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_88 = 7'h58 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_88; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_89 = 7'h59 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_89; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_90 = 7'h5a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_90; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_91 = 7'h5b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_91; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_92 = 7'h5c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_92; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_93 = 7'h5d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_93; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_94 = 7'h5e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_94; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_95 = 7'h5f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_95; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_96 = 7'h60 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_96; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_97 = 7'h61 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_97; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_98 = 7'h62 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_98; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_99 = 7'h63 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_99; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_100 = 7'h64 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_100; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_101 = 7'h65 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_101; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_102 = 7'h66 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_102; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_103 = 7'h67 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_103; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_104 = 7'h68 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_104; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_105 = 7'h69 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_105; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_106 = 7'h6a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_106; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_107 = 7'h6b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_107; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_108 = 7'h6c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_108; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_109 = 7'h6d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_109; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_110 = 7'h6e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_110; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_111 = 7'h6f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_111; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_112 = 7'h70 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_112; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_113 = 7'h71 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_113; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_114 = 7'h72 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_114; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_115 = 7'h73 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_115; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_116 = 7'h74 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_116; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_117 = 7'h75 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_117; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_118 = 7'h76 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_118; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_119 = 7'h77 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_119; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_120 = 7'h78 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_120; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_121 = 7'h79 == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_121; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_122 = 7'h7a == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_122; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_123 = 7'h7b == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_123; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_124 = 7'h7c == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_124; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_125 = 7'h7d == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_125; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_126 = 7'h7e == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_126; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_127 = 7'h7f == io_wrAddr_0[6:0] ? 2'h0 : lvtReg_127; // @[LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 32:28 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_128 = io_wrEna_0 ? _GEN_0 : lvtReg_0; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_129 = io_wrEna_0 ? _GEN_1 : lvtReg_1; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_130 = io_wrEna_0 ? _GEN_2 : lvtReg_2; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_131 = io_wrEna_0 ? _GEN_3 : lvtReg_3; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_132 = io_wrEna_0 ? _GEN_4 : lvtReg_4; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_133 = io_wrEna_0 ? _GEN_5 : lvtReg_5; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_134 = io_wrEna_0 ? _GEN_6 : lvtReg_6; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_135 = io_wrEna_0 ? _GEN_7 : lvtReg_7; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_136 = io_wrEna_0 ? _GEN_8 : lvtReg_8; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_137 = io_wrEna_0 ? _GEN_9 : lvtReg_9; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_138 = io_wrEna_0 ? _GEN_10 : lvtReg_10; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_139 = io_wrEna_0 ? _GEN_11 : lvtReg_11; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_140 = io_wrEna_0 ? _GEN_12 : lvtReg_12; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_141 = io_wrEna_0 ? _GEN_13 : lvtReg_13; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_142 = io_wrEna_0 ? _GEN_14 : lvtReg_14; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_143 = io_wrEna_0 ? _GEN_15 : lvtReg_15; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_144 = io_wrEna_0 ? _GEN_16 : lvtReg_16; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_145 = io_wrEna_0 ? _GEN_17 : lvtReg_17; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_146 = io_wrEna_0 ? _GEN_18 : lvtReg_18; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_147 = io_wrEna_0 ? _GEN_19 : lvtReg_19; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_148 = io_wrEna_0 ? _GEN_20 : lvtReg_20; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_149 = io_wrEna_0 ? _GEN_21 : lvtReg_21; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_150 = io_wrEna_0 ? _GEN_22 : lvtReg_22; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_151 = io_wrEna_0 ? _GEN_23 : lvtReg_23; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_152 = io_wrEna_0 ? _GEN_24 : lvtReg_24; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_153 = io_wrEna_0 ? _GEN_25 : lvtReg_25; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_154 = io_wrEna_0 ? _GEN_26 : lvtReg_26; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_155 = io_wrEna_0 ? _GEN_27 : lvtReg_27; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_156 = io_wrEna_0 ? _GEN_28 : lvtReg_28; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_157 = io_wrEna_0 ? _GEN_29 : lvtReg_29; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_158 = io_wrEna_0 ? _GEN_30 : lvtReg_30; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_159 = io_wrEna_0 ? _GEN_31 : lvtReg_31; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_160 = io_wrEna_0 ? _GEN_32 : lvtReg_32; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_161 = io_wrEna_0 ? _GEN_33 : lvtReg_33; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_162 = io_wrEna_0 ? _GEN_34 : lvtReg_34; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_163 = io_wrEna_0 ? _GEN_35 : lvtReg_35; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_164 = io_wrEna_0 ? _GEN_36 : lvtReg_36; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_165 = io_wrEna_0 ? _GEN_37 : lvtReg_37; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_166 = io_wrEna_0 ? _GEN_38 : lvtReg_38; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_167 = io_wrEna_0 ? _GEN_39 : lvtReg_39; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_168 = io_wrEna_0 ? _GEN_40 : lvtReg_40; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_169 = io_wrEna_0 ? _GEN_41 : lvtReg_41; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_170 = io_wrEna_0 ? _GEN_42 : lvtReg_42; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_171 = io_wrEna_0 ? _GEN_43 : lvtReg_43; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_172 = io_wrEna_0 ? _GEN_44 : lvtReg_44; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_173 = io_wrEna_0 ? _GEN_45 : lvtReg_45; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_174 = io_wrEna_0 ? _GEN_46 : lvtReg_46; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_175 = io_wrEna_0 ? _GEN_47 : lvtReg_47; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_176 = io_wrEna_0 ? _GEN_48 : lvtReg_48; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_177 = io_wrEna_0 ? _GEN_49 : lvtReg_49; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_178 = io_wrEna_0 ? _GEN_50 : lvtReg_50; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_179 = io_wrEna_0 ? _GEN_51 : lvtReg_51; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_180 = io_wrEna_0 ? _GEN_52 : lvtReg_52; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_181 = io_wrEna_0 ? _GEN_53 : lvtReg_53; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_182 = io_wrEna_0 ? _GEN_54 : lvtReg_54; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_183 = io_wrEna_0 ? _GEN_55 : lvtReg_55; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_184 = io_wrEna_0 ? _GEN_56 : lvtReg_56; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_185 = io_wrEna_0 ? _GEN_57 : lvtReg_57; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_186 = io_wrEna_0 ? _GEN_58 : lvtReg_58; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_187 = io_wrEna_0 ? _GEN_59 : lvtReg_59; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_188 = io_wrEna_0 ? _GEN_60 : lvtReg_60; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_189 = io_wrEna_0 ? _GEN_61 : lvtReg_61; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_190 = io_wrEna_0 ? _GEN_62 : lvtReg_62; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_191 = io_wrEna_0 ? _GEN_63 : lvtReg_63; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_192 = io_wrEna_0 ? _GEN_64 : lvtReg_64; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_193 = io_wrEna_0 ? _GEN_65 : lvtReg_65; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_194 = io_wrEna_0 ? _GEN_66 : lvtReg_66; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_195 = io_wrEna_0 ? _GEN_67 : lvtReg_67; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_196 = io_wrEna_0 ? _GEN_68 : lvtReg_68; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_197 = io_wrEna_0 ? _GEN_69 : lvtReg_69; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_198 = io_wrEna_0 ? _GEN_70 : lvtReg_70; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_199 = io_wrEna_0 ? _GEN_71 : lvtReg_71; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_200 = io_wrEna_0 ? _GEN_72 : lvtReg_72; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_201 = io_wrEna_0 ? _GEN_73 : lvtReg_73; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_202 = io_wrEna_0 ? _GEN_74 : lvtReg_74; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_203 = io_wrEna_0 ? _GEN_75 : lvtReg_75; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_204 = io_wrEna_0 ? _GEN_76 : lvtReg_76; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_205 = io_wrEna_0 ? _GEN_77 : lvtReg_77; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_206 = io_wrEna_0 ? _GEN_78 : lvtReg_78; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_207 = io_wrEna_0 ? _GEN_79 : lvtReg_79; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_208 = io_wrEna_0 ? _GEN_80 : lvtReg_80; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_209 = io_wrEna_0 ? _GEN_81 : lvtReg_81; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_210 = io_wrEna_0 ? _GEN_82 : lvtReg_82; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_211 = io_wrEna_0 ? _GEN_83 : lvtReg_83; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_212 = io_wrEna_0 ? _GEN_84 : lvtReg_84; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_213 = io_wrEna_0 ? _GEN_85 : lvtReg_85; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_214 = io_wrEna_0 ? _GEN_86 : lvtReg_86; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_215 = io_wrEna_0 ? _GEN_87 : lvtReg_87; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_216 = io_wrEna_0 ? _GEN_88 : lvtReg_88; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_217 = io_wrEna_0 ? _GEN_89 : lvtReg_89; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_218 = io_wrEna_0 ? _GEN_90 : lvtReg_90; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_219 = io_wrEna_0 ? _GEN_91 : lvtReg_91; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_220 = io_wrEna_0 ? _GEN_92 : lvtReg_92; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_221 = io_wrEna_0 ? _GEN_93 : lvtReg_93; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_222 = io_wrEna_0 ? _GEN_94 : lvtReg_94; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_223 = io_wrEna_0 ? _GEN_95 : lvtReg_95; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_224 = io_wrEna_0 ? _GEN_96 : lvtReg_96; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_225 = io_wrEna_0 ? _GEN_97 : lvtReg_97; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_226 = io_wrEna_0 ? _GEN_98 : lvtReg_98; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_227 = io_wrEna_0 ? _GEN_99 : lvtReg_99; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_228 = io_wrEna_0 ? _GEN_100 : lvtReg_100; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_229 = io_wrEna_0 ? _GEN_101 : lvtReg_101; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_230 = io_wrEna_0 ? _GEN_102 : lvtReg_102; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_231 = io_wrEna_0 ? _GEN_103 : lvtReg_103; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_232 = io_wrEna_0 ? _GEN_104 : lvtReg_104; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_233 = io_wrEna_0 ? _GEN_105 : lvtReg_105; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_234 = io_wrEna_0 ? _GEN_106 : lvtReg_106; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_235 = io_wrEna_0 ? _GEN_107 : lvtReg_107; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_236 = io_wrEna_0 ? _GEN_108 : lvtReg_108; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_237 = io_wrEna_0 ? _GEN_109 : lvtReg_109; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_238 = io_wrEna_0 ? _GEN_110 : lvtReg_110; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_239 = io_wrEna_0 ? _GEN_111 : lvtReg_111; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_240 = io_wrEna_0 ? _GEN_112 : lvtReg_112; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_241 = io_wrEna_0 ? _GEN_113 : lvtReg_113; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_242 = io_wrEna_0 ? _GEN_114 : lvtReg_114; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_243 = io_wrEna_0 ? _GEN_115 : lvtReg_115; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_244 = io_wrEna_0 ? _GEN_116 : lvtReg_116; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_245 = io_wrEna_0 ? _GEN_117 : lvtReg_117; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_246 = io_wrEna_0 ? _GEN_118 : lvtReg_118; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_247 = io_wrEna_0 ? _GEN_119 : lvtReg_119; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_248 = io_wrEna_0 ? _GEN_120 : lvtReg_120; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_249 = io_wrEna_0 ? _GEN_121 : lvtReg_121; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_250 = io_wrEna_0 ? _GEN_122 : lvtReg_122; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_251 = io_wrEna_0 ? _GEN_123 : lvtReg_123; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_252 = io_wrEna_0 ? _GEN_124 : lvtReg_124; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_253 = io_wrEna_0 ? _GEN_125 : lvtReg_125; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_254 = io_wrEna_0 ? _GEN_126 : lvtReg_126; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_255 = io_wrEna_0 ? _GEN_127 : lvtReg_127; // @[LVTMultiPortRams.scala 31:34 LVTMultiPortRams.scala 28:23]
  wire [1:0] _GEN_513 = 7'h1 == io_rdAddr_0[6:0] ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_514 = 7'h2 == io_rdAddr_0[6:0] ? lvtReg_2 : _GEN_513; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_515 = 7'h3 == io_rdAddr_0[6:0] ? lvtReg_3 : _GEN_514; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_516 = 7'h4 == io_rdAddr_0[6:0] ? lvtReg_4 : _GEN_515; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_517 = 7'h5 == io_rdAddr_0[6:0] ? lvtReg_5 : _GEN_516; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_518 = 7'h6 == io_rdAddr_0[6:0] ? lvtReg_6 : _GEN_517; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_519 = 7'h7 == io_rdAddr_0[6:0] ? lvtReg_7 : _GEN_518; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_520 = 7'h8 == io_rdAddr_0[6:0] ? lvtReg_8 : _GEN_519; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_521 = 7'h9 == io_rdAddr_0[6:0] ? lvtReg_9 : _GEN_520; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_522 = 7'ha == io_rdAddr_0[6:0] ? lvtReg_10 : _GEN_521; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_523 = 7'hb == io_rdAddr_0[6:0] ? lvtReg_11 : _GEN_522; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_524 = 7'hc == io_rdAddr_0[6:0] ? lvtReg_12 : _GEN_523; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_525 = 7'hd == io_rdAddr_0[6:0] ? lvtReg_13 : _GEN_524; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_526 = 7'he == io_rdAddr_0[6:0] ? lvtReg_14 : _GEN_525; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_527 = 7'hf == io_rdAddr_0[6:0] ? lvtReg_15 : _GEN_526; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_528 = 7'h10 == io_rdAddr_0[6:0] ? lvtReg_16 : _GEN_527; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_529 = 7'h11 == io_rdAddr_0[6:0] ? lvtReg_17 : _GEN_528; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_530 = 7'h12 == io_rdAddr_0[6:0] ? lvtReg_18 : _GEN_529; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_531 = 7'h13 == io_rdAddr_0[6:0] ? lvtReg_19 : _GEN_530; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_532 = 7'h14 == io_rdAddr_0[6:0] ? lvtReg_20 : _GEN_531; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_533 = 7'h15 == io_rdAddr_0[6:0] ? lvtReg_21 : _GEN_532; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_534 = 7'h16 == io_rdAddr_0[6:0] ? lvtReg_22 : _GEN_533; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_535 = 7'h17 == io_rdAddr_0[6:0] ? lvtReg_23 : _GEN_534; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_536 = 7'h18 == io_rdAddr_0[6:0] ? lvtReg_24 : _GEN_535; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_537 = 7'h19 == io_rdAddr_0[6:0] ? lvtReg_25 : _GEN_536; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_538 = 7'h1a == io_rdAddr_0[6:0] ? lvtReg_26 : _GEN_537; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_539 = 7'h1b == io_rdAddr_0[6:0] ? lvtReg_27 : _GEN_538; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_540 = 7'h1c == io_rdAddr_0[6:0] ? lvtReg_28 : _GEN_539; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_541 = 7'h1d == io_rdAddr_0[6:0] ? lvtReg_29 : _GEN_540; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_542 = 7'h1e == io_rdAddr_0[6:0] ? lvtReg_30 : _GEN_541; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_543 = 7'h1f == io_rdAddr_0[6:0] ? lvtReg_31 : _GEN_542; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_544 = 7'h20 == io_rdAddr_0[6:0] ? lvtReg_32 : _GEN_543; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_545 = 7'h21 == io_rdAddr_0[6:0] ? lvtReg_33 : _GEN_544; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_546 = 7'h22 == io_rdAddr_0[6:0] ? lvtReg_34 : _GEN_545; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_547 = 7'h23 == io_rdAddr_0[6:0] ? lvtReg_35 : _GEN_546; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_548 = 7'h24 == io_rdAddr_0[6:0] ? lvtReg_36 : _GEN_547; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_549 = 7'h25 == io_rdAddr_0[6:0] ? lvtReg_37 : _GEN_548; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_550 = 7'h26 == io_rdAddr_0[6:0] ? lvtReg_38 : _GEN_549; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_551 = 7'h27 == io_rdAddr_0[6:0] ? lvtReg_39 : _GEN_550; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_552 = 7'h28 == io_rdAddr_0[6:0] ? lvtReg_40 : _GEN_551; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_553 = 7'h29 == io_rdAddr_0[6:0] ? lvtReg_41 : _GEN_552; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_554 = 7'h2a == io_rdAddr_0[6:0] ? lvtReg_42 : _GEN_553; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_555 = 7'h2b == io_rdAddr_0[6:0] ? lvtReg_43 : _GEN_554; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_556 = 7'h2c == io_rdAddr_0[6:0] ? lvtReg_44 : _GEN_555; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_557 = 7'h2d == io_rdAddr_0[6:0] ? lvtReg_45 : _GEN_556; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_558 = 7'h2e == io_rdAddr_0[6:0] ? lvtReg_46 : _GEN_557; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_559 = 7'h2f == io_rdAddr_0[6:0] ? lvtReg_47 : _GEN_558; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_560 = 7'h30 == io_rdAddr_0[6:0] ? lvtReg_48 : _GEN_559; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_561 = 7'h31 == io_rdAddr_0[6:0] ? lvtReg_49 : _GEN_560; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_562 = 7'h32 == io_rdAddr_0[6:0] ? lvtReg_50 : _GEN_561; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_563 = 7'h33 == io_rdAddr_0[6:0] ? lvtReg_51 : _GEN_562; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_564 = 7'h34 == io_rdAddr_0[6:0] ? lvtReg_52 : _GEN_563; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_565 = 7'h35 == io_rdAddr_0[6:0] ? lvtReg_53 : _GEN_564; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_566 = 7'h36 == io_rdAddr_0[6:0] ? lvtReg_54 : _GEN_565; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_567 = 7'h37 == io_rdAddr_0[6:0] ? lvtReg_55 : _GEN_566; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_568 = 7'h38 == io_rdAddr_0[6:0] ? lvtReg_56 : _GEN_567; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_569 = 7'h39 == io_rdAddr_0[6:0] ? lvtReg_57 : _GEN_568; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_570 = 7'h3a == io_rdAddr_0[6:0] ? lvtReg_58 : _GEN_569; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_571 = 7'h3b == io_rdAddr_0[6:0] ? lvtReg_59 : _GEN_570; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_572 = 7'h3c == io_rdAddr_0[6:0] ? lvtReg_60 : _GEN_571; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_573 = 7'h3d == io_rdAddr_0[6:0] ? lvtReg_61 : _GEN_572; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_574 = 7'h3e == io_rdAddr_0[6:0] ? lvtReg_62 : _GEN_573; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_575 = 7'h3f == io_rdAddr_0[6:0] ? lvtReg_63 : _GEN_574; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_576 = 7'h40 == io_rdAddr_0[6:0] ? lvtReg_64 : _GEN_575; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_577 = 7'h41 == io_rdAddr_0[6:0] ? lvtReg_65 : _GEN_576; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_578 = 7'h42 == io_rdAddr_0[6:0] ? lvtReg_66 : _GEN_577; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_579 = 7'h43 == io_rdAddr_0[6:0] ? lvtReg_67 : _GEN_578; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_580 = 7'h44 == io_rdAddr_0[6:0] ? lvtReg_68 : _GEN_579; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_581 = 7'h45 == io_rdAddr_0[6:0] ? lvtReg_69 : _GEN_580; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_582 = 7'h46 == io_rdAddr_0[6:0] ? lvtReg_70 : _GEN_581; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_583 = 7'h47 == io_rdAddr_0[6:0] ? lvtReg_71 : _GEN_582; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_584 = 7'h48 == io_rdAddr_0[6:0] ? lvtReg_72 : _GEN_583; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_585 = 7'h49 == io_rdAddr_0[6:0] ? lvtReg_73 : _GEN_584; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_586 = 7'h4a == io_rdAddr_0[6:0] ? lvtReg_74 : _GEN_585; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_587 = 7'h4b == io_rdAddr_0[6:0] ? lvtReg_75 : _GEN_586; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_588 = 7'h4c == io_rdAddr_0[6:0] ? lvtReg_76 : _GEN_587; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_589 = 7'h4d == io_rdAddr_0[6:0] ? lvtReg_77 : _GEN_588; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_590 = 7'h4e == io_rdAddr_0[6:0] ? lvtReg_78 : _GEN_589; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_591 = 7'h4f == io_rdAddr_0[6:0] ? lvtReg_79 : _GEN_590; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_592 = 7'h50 == io_rdAddr_0[6:0] ? lvtReg_80 : _GEN_591; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_593 = 7'h51 == io_rdAddr_0[6:0] ? lvtReg_81 : _GEN_592; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_594 = 7'h52 == io_rdAddr_0[6:0] ? lvtReg_82 : _GEN_593; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_595 = 7'h53 == io_rdAddr_0[6:0] ? lvtReg_83 : _GEN_594; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_596 = 7'h54 == io_rdAddr_0[6:0] ? lvtReg_84 : _GEN_595; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_597 = 7'h55 == io_rdAddr_0[6:0] ? lvtReg_85 : _GEN_596; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_598 = 7'h56 == io_rdAddr_0[6:0] ? lvtReg_86 : _GEN_597; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_599 = 7'h57 == io_rdAddr_0[6:0] ? lvtReg_87 : _GEN_598; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_600 = 7'h58 == io_rdAddr_0[6:0] ? lvtReg_88 : _GEN_599; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_601 = 7'h59 == io_rdAddr_0[6:0] ? lvtReg_89 : _GEN_600; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_602 = 7'h5a == io_rdAddr_0[6:0] ? lvtReg_90 : _GEN_601; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_603 = 7'h5b == io_rdAddr_0[6:0] ? lvtReg_91 : _GEN_602; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_604 = 7'h5c == io_rdAddr_0[6:0] ? lvtReg_92 : _GEN_603; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_605 = 7'h5d == io_rdAddr_0[6:0] ? lvtReg_93 : _GEN_604; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_606 = 7'h5e == io_rdAddr_0[6:0] ? lvtReg_94 : _GEN_605; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_607 = 7'h5f == io_rdAddr_0[6:0] ? lvtReg_95 : _GEN_606; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_608 = 7'h60 == io_rdAddr_0[6:0] ? lvtReg_96 : _GEN_607; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_609 = 7'h61 == io_rdAddr_0[6:0] ? lvtReg_97 : _GEN_608; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_610 = 7'h62 == io_rdAddr_0[6:0] ? lvtReg_98 : _GEN_609; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_611 = 7'h63 == io_rdAddr_0[6:0] ? lvtReg_99 : _GEN_610; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_612 = 7'h64 == io_rdAddr_0[6:0] ? lvtReg_100 : _GEN_611; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_613 = 7'h65 == io_rdAddr_0[6:0] ? lvtReg_101 : _GEN_612; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_614 = 7'h66 == io_rdAddr_0[6:0] ? lvtReg_102 : _GEN_613; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_615 = 7'h67 == io_rdAddr_0[6:0] ? lvtReg_103 : _GEN_614; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_616 = 7'h68 == io_rdAddr_0[6:0] ? lvtReg_104 : _GEN_615; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_617 = 7'h69 == io_rdAddr_0[6:0] ? lvtReg_105 : _GEN_616; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_618 = 7'h6a == io_rdAddr_0[6:0] ? lvtReg_106 : _GEN_617; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_619 = 7'h6b == io_rdAddr_0[6:0] ? lvtReg_107 : _GEN_618; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_620 = 7'h6c == io_rdAddr_0[6:0] ? lvtReg_108 : _GEN_619; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_621 = 7'h6d == io_rdAddr_0[6:0] ? lvtReg_109 : _GEN_620; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_622 = 7'h6e == io_rdAddr_0[6:0] ? lvtReg_110 : _GEN_621; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_623 = 7'h6f == io_rdAddr_0[6:0] ? lvtReg_111 : _GEN_622; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_624 = 7'h70 == io_rdAddr_0[6:0] ? lvtReg_112 : _GEN_623; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_625 = 7'h71 == io_rdAddr_0[6:0] ? lvtReg_113 : _GEN_624; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_626 = 7'h72 == io_rdAddr_0[6:0] ? lvtReg_114 : _GEN_625; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_627 = 7'h73 == io_rdAddr_0[6:0] ? lvtReg_115 : _GEN_626; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_628 = 7'h74 == io_rdAddr_0[6:0] ? lvtReg_116 : _GEN_627; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_629 = 7'h75 == io_rdAddr_0[6:0] ? lvtReg_117 : _GEN_628; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_630 = 7'h76 == io_rdAddr_0[6:0] ? lvtReg_118 : _GEN_629; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_631 = 7'h77 == io_rdAddr_0[6:0] ? lvtReg_119 : _GEN_630; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_632 = 7'h78 == io_rdAddr_0[6:0] ? lvtReg_120 : _GEN_631; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_633 = 7'h79 == io_rdAddr_0[6:0] ? lvtReg_121 : _GEN_632; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_634 = 7'h7a == io_rdAddr_0[6:0] ? lvtReg_122 : _GEN_633; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_635 = 7'h7b == io_rdAddr_0[6:0] ? lvtReg_123 : _GEN_634; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_636 = 7'h7c == io_rdAddr_0[6:0] ? lvtReg_124 : _GEN_635; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_637 = 7'h7d == io_rdAddr_0[6:0] ? lvtReg_125 : _GEN_636; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_638 = 7'h7e == io_rdAddr_0[6:0] ? lvtReg_126 : _GEN_637; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_641 = 7'h1 == io_rdAddr_1[6:0] ? lvtReg_1 : lvtReg_0; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_642 = 7'h2 == io_rdAddr_1[6:0] ? lvtReg_2 : _GEN_641; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_643 = 7'h3 == io_rdAddr_1[6:0] ? lvtReg_3 : _GEN_642; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_644 = 7'h4 == io_rdAddr_1[6:0] ? lvtReg_4 : _GEN_643; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_645 = 7'h5 == io_rdAddr_1[6:0] ? lvtReg_5 : _GEN_644; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_646 = 7'h6 == io_rdAddr_1[6:0] ? lvtReg_6 : _GEN_645; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_647 = 7'h7 == io_rdAddr_1[6:0] ? lvtReg_7 : _GEN_646; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_648 = 7'h8 == io_rdAddr_1[6:0] ? lvtReg_8 : _GEN_647; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_649 = 7'h9 == io_rdAddr_1[6:0] ? lvtReg_9 : _GEN_648; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_650 = 7'ha == io_rdAddr_1[6:0] ? lvtReg_10 : _GEN_649; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_651 = 7'hb == io_rdAddr_1[6:0] ? lvtReg_11 : _GEN_650; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_652 = 7'hc == io_rdAddr_1[6:0] ? lvtReg_12 : _GEN_651; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_653 = 7'hd == io_rdAddr_1[6:0] ? lvtReg_13 : _GEN_652; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_654 = 7'he == io_rdAddr_1[6:0] ? lvtReg_14 : _GEN_653; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_655 = 7'hf == io_rdAddr_1[6:0] ? lvtReg_15 : _GEN_654; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_656 = 7'h10 == io_rdAddr_1[6:0] ? lvtReg_16 : _GEN_655; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_657 = 7'h11 == io_rdAddr_1[6:0] ? lvtReg_17 : _GEN_656; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_658 = 7'h12 == io_rdAddr_1[6:0] ? lvtReg_18 : _GEN_657; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_659 = 7'h13 == io_rdAddr_1[6:0] ? lvtReg_19 : _GEN_658; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_660 = 7'h14 == io_rdAddr_1[6:0] ? lvtReg_20 : _GEN_659; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_661 = 7'h15 == io_rdAddr_1[6:0] ? lvtReg_21 : _GEN_660; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_662 = 7'h16 == io_rdAddr_1[6:0] ? lvtReg_22 : _GEN_661; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_663 = 7'h17 == io_rdAddr_1[6:0] ? lvtReg_23 : _GEN_662; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_664 = 7'h18 == io_rdAddr_1[6:0] ? lvtReg_24 : _GEN_663; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_665 = 7'h19 == io_rdAddr_1[6:0] ? lvtReg_25 : _GEN_664; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_666 = 7'h1a == io_rdAddr_1[6:0] ? lvtReg_26 : _GEN_665; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_667 = 7'h1b == io_rdAddr_1[6:0] ? lvtReg_27 : _GEN_666; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_668 = 7'h1c == io_rdAddr_1[6:0] ? lvtReg_28 : _GEN_667; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_669 = 7'h1d == io_rdAddr_1[6:0] ? lvtReg_29 : _GEN_668; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_670 = 7'h1e == io_rdAddr_1[6:0] ? lvtReg_30 : _GEN_669; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_671 = 7'h1f == io_rdAddr_1[6:0] ? lvtReg_31 : _GEN_670; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_672 = 7'h20 == io_rdAddr_1[6:0] ? lvtReg_32 : _GEN_671; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_673 = 7'h21 == io_rdAddr_1[6:0] ? lvtReg_33 : _GEN_672; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_674 = 7'h22 == io_rdAddr_1[6:0] ? lvtReg_34 : _GEN_673; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_675 = 7'h23 == io_rdAddr_1[6:0] ? lvtReg_35 : _GEN_674; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_676 = 7'h24 == io_rdAddr_1[6:0] ? lvtReg_36 : _GEN_675; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_677 = 7'h25 == io_rdAddr_1[6:0] ? lvtReg_37 : _GEN_676; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_678 = 7'h26 == io_rdAddr_1[6:0] ? lvtReg_38 : _GEN_677; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_679 = 7'h27 == io_rdAddr_1[6:0] ? lvtReg_39 : _GEN_678; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_680 = 7'h28 == io_rdAddr_1[6:0] ? lvtReg_40 : _GEN_679; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_681 = 7'h29 == io_rdAddr_1[6:0] ? lvtReg_41 : _GEN_680; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_682 = 7'h2a == io_rdAddr_1[6:0] ? lvtReg_42 : _GEN_681; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_683 = 7'h2b == io_rdAddr_1[6:0] ? lvtReg_43 : _GEN_682; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_684 = 7'h2c == io_rdAddr_1[6:0] ? lvtReg_44 : _GEN_683; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_685 = 7'h2d == io_rdAddr_1[6:0] ? lvtReg_45 : _GEN_684; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_686 = 7'h2e == io_rdAddr_1[6:0] ? lvtReg_46 : _GEN_685; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_687 = 7'h2f == io_rdAddr_1[6:0] ? lvtReg_47 : _GEN_686; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_688 = 7'h30 == io_rdAddr_1[6:0] ? lvtReg_48 : _GEN_687; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_689 = 7'h31 == io_rdAddr_1[6:0] ? lvtReg_49 : _GEN_688; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_690 = 7'h32 == io_rdAddr_1[6:0] ? lvtReg_50 : _GEN_689; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_691 = 7'h33 == io_rdAddr_1[6:0] ? lvtReg_51 : _GEN_690; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_692 = 7'h34 == io_rdAddr_1[6:0] ? lvtReg_52 : _GEN_691; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_693 = 7'h35 == io_rdAddr_1[6:0] ? lvtReg_53 : _GEN_692; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_694 = 7'h36 == io_rdAddr_1[6:0] ? lvtReg_54 : _GEN_693; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_695 = 7'h37 == io_rdAddr_1[6:0] ? lvtReg_55 : _GEN_694; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_696 = 7'h38 == io_rdAddr_1[6:0] ? lvtReg_56 : _GEN_695; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_697 = 7'h39 == io_rdAddr_1[6:0] ? lvtReg_57 : _GEN_696; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_698 = 7'h3a == io_rdAddr_1[6:0] ? lvtReg_58 : _GEN_697; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_699 = 7'h3b == io_rdAddr_1[6:0] ? lvtReg_59 : _GEN_698; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_700 = 7'h3c == io_rdAddr_1[6:0] ? lvtReg_60 : _GEN_699; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_701 = 7'h3d == io_rdAddr_1[6:0] ? lvtReg_61 : _GEN_700; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_702 = 7'h3e == io_rdAddr_1[6:0] ? lvtReg_62 : _GEN_701; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_703 = 7'h3f == io_rdAddr_1[6:0] ? lvtReg_63 : _GEN_702; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_704 = 7'h40 == io_rdAddr_1[6:0] ? lvtReg_64 : _GEN_703; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_705 = 7'h41 == io_rdAddr_1[6:0] ? lvtReg_65 : _GEN_704; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_706 = 7'h42 == io_rdAddr_1[6:0] ? lvtReg_66 : _GEN_705; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_707 = 7'h43 == io_rdAddr_1[6:0] ? lvtReg_67 : _GEN_706; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_708 = 7'h44 == io_rdAddr_1[6:0] ? lvtReg_68 : _GEN_707; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_709 = 7'h45 == io_rdAddr_1[6:0] ? lvtReg_69 : _GEN_708; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_710 = 7'h46 == io_rdAddr_1[6:0] ? lvtReg_70 : _GEN_709; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_711 = 7'h47 == io_rdAddr_1[6:0] ? lvtReg_71 : _GEN_710; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_712 = 7'h48 == io_rdAddr_1[6:0] ? lvtReg_72 : _GEN_711; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_713 = 7'h49 == io_rdAddr_1[6:0] ? lvtReg_73 : _GEN_712; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_714 = 7'h4a == io_rdAddr_1[6:0] ? lvtReg_74 : _GEN_713; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_715 = 7'h4b == io_rdAddr_1[6:0] ? lvtReg_75 : _GEN_714; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_716 = 7'h4c == io_rdAddr_1[6:0] ? lvtReg_76 : _GEN_715; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_717 = 7'h4d == io_rdAddr_1[6:0] ? lvtReg_77 : _GEN_716; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_718 = 7'h4e == io_rdAddr_1[6:0] ? lvtReg_78 : _GEN_717; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_719 = 7'h4f == io_rdAddr_1[6:0] ? lvtReg_79 : _GEN_718; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_720 = 7'h50 == io_rdAddr_1[6:0] ? lvtReg_80 : _GEN_719; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_721 = 7'h51 == io_rdAddr_1[6:0] ? lvtReg_81 : _GEN_720; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_722 = 7'h52 == io_rdAddr_1[6:0] ? lvtReg_82 : _GEN_721; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_723 = 7'h53 == io_rdAddr_1[6:0] ? lvtReg_83 : _GEN_722; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_724 = 7'h54 == io_rdAddr_1[6:0] ? lvtReg_84 : _GEN_723; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_725 = 7'h55 == io_rdAddr_1[6:0] ? lvtReg_85 : _GEN_724; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_726 = 7'h56 == io_rdAddr_1[6:0] ? lvtReg_86 : _GEN_725; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_727 = 7'h57 == io_rdAddr_1[6:0] ? lvtReg_87 : _GEN_726; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_728 = 7'h58 == io_rdAddr_1[6:0] ? lvtReg_88 : _GEN_727; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_729 = 7'h59 == io_rdAddr_1[6:0] ? lvtReg_89 : _GEN_728; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_730 = 7'h5a == io_rdAddr_1[6:0] ? lvtReg_90 : _GEN_729; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_731 = 7'h5b == io_rdAddr_1[6:0] ? lvtReg_91 : _GEN_730; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_732 = 7'h5c == io_rdAddr_1[6:0] ? lvtReg_92 : _GEN_731; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_733 = 7'h5d == io_rdAddr_1[6:0] ? lvtReg_93 : _GEN_732; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_734 = 7'h5e == io_rdAddr_1[6:0] ? lvtReg_94 : _GEN_733; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_735 = 7'h5f == io_rdAddr_1[6:0] ? lvtReg_95 : _GEN_734; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_736 = 7'h60 == io_rdAddr_1[6:0] ? lvtReg_96 : _GEN_735; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_737 = 7'h61 == io_rdAddr_1[6:0] ? lvtReg_97 : _GEN_736; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_738 = 7'h62 == io_rdAddr_1[6:0] ? lvtReg_98 : _GEN_737; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_739 = 7'h63 == io_rdAddr_1[6:0] ? lvtReg_99 : _GEN_738; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_740 = 7'h64 == io_rdAddr_1[6:0] ? lvtReg_100 : _GEN_739; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_741 = 7'h65 == io_rdAddr_1[6:0] ? lvtReg_101 : _GEN_740; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_742 = 7'h66 == io_rdAddr_1[6:0] ? lvtReg_102 : _GEN_741; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_743 = 7'h67 == io_rdAddr_1[6:0] ? lvtReg_103 : _GEN_742; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_744 = 7'h68 == io_rdAddr_1[6:0] ? lvtReg_104 : _GEN_743; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_745 = 7'h69 == io_rdAddr_1[6:0] ? lvtReg_105 : _GEN_744; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_746 = 7'h6a == io_rdAddr_1[6:0] ? lvtReg_106 : _GEN_745; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_747 = 7'h6b == io_rdAddr_1[6:0] ? lvtReg_107 : _GEN_746; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_748 = 7'h6c == io_rdAddr_1[6:0] ? lvtReg_108 : _GEN_747; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_749 = 7'h6d == io_rdAddr_1[6:0] ? lvtReg_109 : _GEN_748; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_750 = 7'h6e == io_rdAddr_1[6:0] ? lvtReg_110 : _GEN_749; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_751 = 7'h6f == io_rdAddr_1[6:0] ? lvtReg_111 : _GEN_750; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_752 = 7'h70 == io_rdAddr_1[6:0] ? lvtReg_112 : _GEN_751; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_753 = 7'h71 == io_rdAddr_1[6:0] ? lvtReg_113 : _GEN_752; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_754 = 7'h72 == io_rdAddr_1[6:0] ? lvtReg_114 : _GEN_753; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_755 = 7'h73 == io_rdAddr_1[6:0] ? lvtReg_115 : _GEN_754; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_756 = 7'h74 == io_rdAddr_1[6:0] ? lvtReg_116 : _GEN_755; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_757 = 7'h75 == io_rdAddr_1[6:0] ? lvtReg_117 : _GEN_756; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_758 = 7'h76 == io_rdAddr_1[6:0] ? lvtReg_118 : _GEN_757; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_759 = 7'h77 == io_rdAddr_1[6:0] ? lvtReg_119 : _GEN_758; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_760 = 7'h78 == io_rdAddr_1[6:0] ? lvtReg_120 : _GEN_759; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_761 = 7'h79 == io_rdAddr_1[6:0] ? lvtReg_121 : _GEN_760; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_762 = 7'h7a == io_rdAddr_1[6:0] ? lvtReg_122 : _GEN_761; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_763 = 7'h7b == io_rdAddr_1[6:0] ? lvtReg_123 : _GEN_762; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_764 = 7'h7c == io_rdAddr_1[6:0] ? lvtReg_124 : _GEN_763; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_765 = 7'h7d == io_rdAddr_1[6:0] ? lvtReg_125 : _GEN_764; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  wire [1:0] _GEN_766 = 7'h7e == io_rdAddr_1[6:0] ? lvtReg_126 : _GEN_765; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_0 = 7'h7f == io_rdAddr_0[6:0] ? lvtReg_127 : _GEN_638; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  assign io_rdIdx_1 = 7'h7f == io_rdAddr_1[6:0] ? lvtReg_127 : _GEN_766; // @[LVTMultiPortRams.scala 37:17 LVTMultiPortRams.scala 37:17]
  always @(posedge clock) begin
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_0 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h0 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_0 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_0 <= _GEN_128;
      end
    end else begin
      lvtReg_0 <= _GEN_128;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_1 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_1 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_1 <= _GEN_129;
      end
    end else begin
      lvtReg_1 <= _GEN_129;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_2 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_2 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_2 <= _GEN_130;
      end
    end else begin
      lvtReg_2 <= _GEN_130;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_3 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_3 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_3 <= _GEN_131;
      end
    end else begin
      lvtReg_3 <= _GEN_131;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_4 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_4 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_4 <= _GEN_132;
      end
    end else begin
      lvtReg_4 <= _GEN_132;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_5 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_5 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_5 <= _GEN_133;
      end
    end else begin
      lvtReg_5 <= _GEN_133;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_6 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_6 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_6 <= _GEN_134;
      end
    end else begin
      lvtReg_6 <= _GEN_134;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_7 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_7 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_7 <= _GEN_135;
      end
    end else begin
      lvtReg_7 <= _GEN_135;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_8 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h8 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_8 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_8 <= _GEN_136;
      end
    end else begin
      lvtReg_8 <= _GEN_136;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_9 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h9 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_9 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_9 <= _GEN_137;
      end
    end else begin
      lvtReg_9 <= _GEN_137;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_10 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'ha == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_10 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_10 <= _GEN_138;
      end
    end else begin
      lvtReg_10 <= _GEN_138;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_11 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'hb == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_11 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_11 <= _GEN_139;
      end
    end else begin
      lvtReg_11 <= _GEN_139;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_12 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'hc == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_12 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_12 <= _GEN_140;
      end
    end else begin
      lvtReg_12 <= _GEN_140;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_13 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'hd == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_13 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_13 <= _GEN_141;
      end
    end else begin
      lvtReg_13 <= _GEN_141;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_14 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'he == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_14 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_14 <= _GEN_142;
      end
    end else begin
      lvtReg_14 <= _GEN_142;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_15 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'hf == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_15 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_15 <= _GEN_143;
      end
    end else begin
      lvtReg_15 <= _GEN_143;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_16 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h10 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_16 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_16 <= _GEN_144;
      end
    end else begin
      lvtReg_16 <= _GEN_144;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_17 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h11 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_17 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_17 <= _GEN_145;
      end
    end else begin
      lvtReg_17 <= _GEN_145;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_18 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h12 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_18 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_18 <= _GEN_146;
      end
    end else begin
      lvtReg_18 <= _GEN_146;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_19 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h13 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_19 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_19 <= _GEN_147;
      end
    end else begin
      lvtReg_19 <= _GEN_147;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_20 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h14 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_20 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_20 <= _GEN_148;
      end
    end else begin
      lvtReg_20 <= _GEN_148;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_21 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h15 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_21 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_21 <= _GEN_149;
      end
    end else begin
      lvtReg_21 <= _GEN_149;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_22 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h16 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_22 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_22 <= _GEN_150;
      end
    end else begin
      lvtReg_22 <= _GEN_150;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_23 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h17 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_23 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_23 <= _GEN_151;
      end
    end else begin
      lvtReg_23 <= _GEN_151;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_24 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h18 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_24 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_24 <= _GEN_152;
      end
    end else begin
      lvtReg_24 <= _GEN_152;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_25 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h19 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_25 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_25 <= _GEN_153;
      end
    end else begin
      lvtReg_25 <= _GEN_153;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_26 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_26 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_26 <= _GEN_154;
      end
    end else begin
      lvtReg_26 <= _GEN_154;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_27 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_27 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_27 <= _GEN_155;
      end
    end else begin
      lvtReg_27 <= _GEN_155;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_28 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_28 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_28 <= _GEN_156;
      end
    end else begin
      lvtReg_28 <= _GEN_156;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_29 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_29 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_29 <= _GEN_157;
      end
    end else begin
      lvtReg_29 <= _GEN_157;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_30 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_30 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_30 <= _GEN_158;
      end
    end else begin
      lvtReg_30 <= _GEN_158;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_31 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h1f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_31 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_31 <= _GEN_159;
      end
    end else begin
      lvtReg_31 <= _GEN_159;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_32 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h20 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_32 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_32 <= _GEN_160;
      end
    end else begin
      lvtReg_32 <= _GEN_160;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_33 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h21 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_33 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_33 <= _GEN_161;
      end
    end else begin
      lvtReg_33 <= _GEN_161;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_34 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h22 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_34 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_34 <= _GEN_162;
      end
    end else begin
      lvtReg_34 <= _GEN_162;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_35 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h23 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_35 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_35 <= _GEN_163;
      end
    end else begin
      lvtReg_35 <= _GEN_163;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_36 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h24 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_36 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_36 <= _GEN_164;
      end
    end else begin
      lvtReg_36 <= _GEN_164;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_37 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h25 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_37 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_37 <= _GEN_165;
      end
    end else begin
      lvtReg_37 <= _GEN_165;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_38 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h26 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_38 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_38 <= _GEN_166;
      end
    end else begin
      lvtReg_38 <= _GEN_166;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_39 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h27 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_39 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_39 <= _GEN_167;
      end
    end else begin
      lvtReg_39 <= _GEN_167;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_40 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h28 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_40 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_40 <= _GEN_168;
      end
    end else begin
      lvtReg_40 <= _GEN_168;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_41 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h29 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_41 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_41 <= _GEN_169;
      end
    end else begin
      lvtReg_41 <= _GEN_169;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_42 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_42 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_42 <= _GEN_170;
      end
    end else begin
      lvtReg_42 <= _GEN_170;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_43 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_43 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_43 <= _GEN_171;
      end
    end else begin
      lvtReg_43 <= _GEN_171;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_44 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_44 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_44 <= _GEN_172;
      end
    end else begin
      lvtReg_44 <= _GEN_172;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_45 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_45 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_45 <= _GEN_173;
      end
    end else begin
      lvtReg_45 <= _GEN_173;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_46 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_46 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_46 <= _GEN_174;
      end
    end else begin
      lvtReg_46 <= _GEN_174;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_47 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h2f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_47 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_47 <= _GEN_175;
      end
    end else begin
      lvtReg_47 <= _GEN_175;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_48 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h30 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_48 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_48 <= _GEN_176;
      end
    end else begin
      lvtReg_48 <= _GEN_176;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_49 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h31 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_49 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_49 <= _GEN_177;
      end
    end else begin
      lvtReg_49 <= _GEN_177;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_50 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h32 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_50 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_50 <= _GEN_178;
      end
    end else begin
      lvtReg_50 <= _GEN_178;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_51 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h33 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_51 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_51 <= _GEN_179;
      end
    end else begin
      lvtReg_51 <= _GEN_179;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_52 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h34 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_52 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_52 <= _GEN_180;
      end
    end else begin
      lvtReg_52 <= _GEN_180;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_53 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h35 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_53 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_53 <= _GEN_181;
      end
    end else begin
      lvtReg_53 <= _GEN_181;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_54 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h36 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_54 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_54 <= _GEN_182;
      end
    end else begin
      lvtReg_54 <= _GEN_182;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_55 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h37 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_55 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_55 <= _GEN_183;
      end
    end else begin
      lvtReg_55 <= _GEN_183;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_56 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h38 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_56 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_56 <= _GEN_184;
      end
    end else begin
      lvtReg_56 <= _GEN_184;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_57 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h39 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_57 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_57 <= _GEN_185;
      end
    end else begin
      lvtReg_57 <= _GEN_185;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_58 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_58 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_58 <= _GEN_186;
      end
    end else begin
      lvtReg_58 <= _GEN_186;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_59 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_59 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_59 <= _GEN_187;
      end
    end else begin
      lvtReg_59 <= _GEN_187;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_60 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_60 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_60 <= _GEN_188;
      end
    end else begin
      lvtReg_60 <= _GEN_188;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_61 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_61 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_61 <= _GEN_189;
      end
    end else begin
      lvtReg_61 <= _GEN_189;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_62 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_62 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_62 <= _GEN_190;
      end
    end else begin
      lvtReg_62 <= _GEN_190;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_63 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h3f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_63 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_63 <= _GEN_191;
      end
    end else begin
      lvtReg_63 <= _GEN_191;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_64 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h40 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_64 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_64 <= _GEN_192;
      end
    end else begin
      lvtReg_64 <= _GEN_192;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_65 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h41 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_65 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_65 <= _GEN_193;
      end
    end else begin
      lvtReg_65 <= _GEN_193;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_66 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h42 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_66 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_66 <= _GEN_194;
      end
    end else begin
      lvtReg_66 <= _GEN_194;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_67 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h43 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_67 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_67 <= _GEN_195;
      end
    end else begin
      lvtReg_67 <= _GEN_195;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_68 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h44 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_68 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_68 <= _GEN_196;
      end
    end else begin
      lvtReg_68 <= _GEN_196;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_69 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h45 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_69 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_69 <= _GEN_197;
      end
    end else begin
      lvtReg_69 <= _GEN_197;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_70 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h46 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_70 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_70 <= _GEN_198;
      end
    end else begin
      lvtReg_70 <= _GEN_198;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_71 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h47 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_71 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_71 <= _GEN_199;
      end
    end else begin
      lvtReg_71 <= _GEN_199;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_72 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h48 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_72 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_72 <= _GEN_200;
      end
    end else begin
      lvtReg_72 <= _GEN_200;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_73 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h49 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_73 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_73 <= _GEN_201;
      end
    end else begin
      lvtReg_73 <= _GEN_201;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_74 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_74 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_74 <= _GEN_202;
      end
    end else begin
      lvtReg_74 <= _GEN_202;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_75 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_75 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_75 <= _GEN_203;
      end
    end else begin
      lvtReg_75 <= _GEN_203;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_76 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_76 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_76 <= _GEN_204;
      end
    end else begin
      lvtReg_76 <= _GEN_204;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_77 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_77 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_77 <= _GEN_205;
      end
    end else begin
      lvtReg_77 <= _GEN_205;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_78 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_78 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_78 <= _GEN_206;
      end
    end else begin
      lvtReg_78 <= _GEN_206;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_79 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h4f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_79 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_79 <= _GEN_207;
      end
    end else begin
      lvtReg_79 <= _GEN_207;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_80 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h50 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_80 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_80 <= _GEN_208;
      end
    end else begin
      lvtReg_80 <= _GEN_208;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_81 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h51 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_81 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_81 <= _GEN_209;
      end
    end else begin
      lvtReg_81 <= _GEN_209;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_82 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h52 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_82 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_82 <= _GEN_210;
      end
    end else begin
      lvtReg_82 <= _GEN_210;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_83 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h53 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_83 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_83 <= _GEN_211;
      end
    end else begin
      lvtReg_83 <= _GEN_211;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_84 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h54 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_84 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_84 <= _GEN_212;
      end
    end else begin
      lvtReg_84 <= _GEN_212;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_85 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h55 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_85 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_85 <= _GEN_213;
      end
    end else begin
      lvtReg_85 <= _GEN_213;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_86 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h56 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_86 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_86 <= _GEN_214;
      end
    end else begin
      lvtReg_86 <= _GEN_214;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_87 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h57 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_87 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_87 <= _GEN_215;
      end
    end else begin
      lvtReg_87 <= _GEN_215;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_88 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h58 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_88 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_88 <= _GEN_216;
      end
    end else begin
      lvtReg_88 <= _GEN_216;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_89 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h59 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_89 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_89 <= _GEN_217;
      end
    end else begin
      lvtReg_89 <= _GEN_217;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_90 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_90 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_90 <= _GEN_218;
      end
    end else begin
      lvtReg_90 <= _GEN_218;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_91 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_91 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_91 <= _GEN_219;
      end
    end else begin
      lvtReg_91 <= _GEN_219;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_92 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_92 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_92 <= _GEN_220;
      end
    end else begin
      lvtReg_92 <= _GEN_220;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_93 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_93 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_93 <= _GEN_221;
      end
    end else begin
      lvtReg_93 <= _GEN_221;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_94 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_94 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_94 <= _GEN_222;
      end
    end else begin
      lvtReg_94 <= _GEN_222;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_95 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h5f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_95 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_95 <= _GEN_223;
      end
    end else begin
      lvtReg_95 <= _GEN_223;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_96 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h60 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_96 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_96 <= _GEN_224;
      end
    end else begin
      lvtReg_96 <= _GEN_224;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_97 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h61 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_97 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_97 <= _GEN_225;
      end
    end else begin
      lvtReg_97 <= _GEN_225;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_98 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h62 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_98 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_98 <= _GEN_226;
      end
    end else begin
      lvtReg_98 <= _GEN_226;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_99 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h63 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_99 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_99 <= _GEN_227;
      end
    end else begin
      lvtReg_99 <= _GEN_227;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_100 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h64 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_100 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_100 <= _GEN_228;
      end
    end else begin
      lvtReg_100 <= _GEN_228;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_101 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h65 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_101 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_101 <= _GEN_229;
      end
    end else begin
      lvtReg_101 <= _GEN_229;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_102 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h66 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_102 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_102 <= _GEN_230;
      end
    end else begin
      lvtReg_102 <= _GEN_230;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_103 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h67 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_103 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_103 <= _GEN_231;
      end
    end else begin
      lvtReg_103 <= _GEN_231;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_104 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h68 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_104 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_104 <= _GEN_232;
      end
    end else begin
      lvtReg_104 <= _GEN_232;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_105 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h69 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_105 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_105 <= _GEN_233;
      end
    end else begin
      lvtReg_105 <= _GEN_233;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_106 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_106 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_106 <= _GEN_234;
      end
    end else begin
      lvtReg_106 <= _GEN_234;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_107 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_107 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_107 <= _GEN_235;
      end
    end else begin
      lvtReg_107 <= _GEN_235;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_108 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_108 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_108 <= _GEN_236;
      end
    end else begin
      lvtReg_108 <= _GEN_236;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_109 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_109 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_109 <= _GEN_237;
      end
    end else begin
      lvtReg_109 <= _GEN_237;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_110 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_110 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_110 <= _GEN_238;
      end
    end else begin
      lvtReg_110 <= _GEN_238;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_111 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h6f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_111 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_111 <= _GEN_239;
      end
    end else begin
      lvtReg_111 <= _GEN_239;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_112 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h70 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_112 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_112 <= _GEN_240;
      end
    end else begin
      lvtReg_112 <= _GEN_240;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_113 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h71 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_113 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_113 <= _GEN_241;
      end
    end else begin
      lvtReg_113 <= _GEN_241;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_114 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h72 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_114 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_114 <= _GEN_242;
      end
    end else begin
      lvtReg_114 <= _GEN_242;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_115 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h73 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_115 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_115 <= _GEN_243;
      end
    end else begin
      lvtReg_115 <= _GEN_243;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_116 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h74 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_116 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_116 <= _GEN_244;
      end
    end else begin
      lvtReg_116 <= _GEN_244;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_117 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h75 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_117 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_117 <= _GEN_245;
      end
    end else begin
      lvtReg_117 <= _GEN_245;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_118 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h76 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_118 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_118 <= _GEN_246;
      end
    end else begin
      lvtReg_118 <= _GEN_246;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_119 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h77 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_119 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_119 <= _GEN_247;
      end
    end else begin
      lvtReg_119 <= _GEN_247;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_120 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h78 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_120 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_120 <= _GEN_248;
      end
    end else begin
      lvtReg_120 <= _GEN_248;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_121 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h79 == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_121 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_121 <= _GEN_249;
      end
    end else begin
      lvtReg_121 <= _GEN_249;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_122 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7a == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_122 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_122 <= _GEN_250;
      end
    end else begin
      lvtReg_122 <= _GEN_250;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_123 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7b == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_123 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_123 <= _GEN_251;
      end
    end else begin
      lvtReg_123 <= _GEN_251;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_124 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7c == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_124 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_124 <= _GEN_252;
      end
    end else begin
      lvtReg_124 <= _GEN_252;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_125 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7d == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_125 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_125 <= _GEN_253;
      end
    end else begin
      lvtReg_125 <= _GEN_253;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_126 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7e == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_126 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_126 <= _GEN_254;
      end
    end else begin
      lvtReg_126 <= _GEN_254;
    end
    if (reset) begin // @[LVTMultiPortRams.scala 28:23]
      lvtReg_127 <= 2'h0; // @[LVTMultiPortRams.scala 28:23]
    end else if (io_wrEna_1) begin // @[LVTMultiPortRams.scala 31:34]
      if (7'h7f == io_wrAddr_1[6:0]) begin // @[LVTMultiPortRams.scala 32:28]
        lvtReg_127 <= 2'h1; // @[LVTMultiPortRams.scala 32:28]
      end else begin
        lvtReg_127 <= _GEN_255;
      end
    end else begin
      lvtReg_127 <= _GEN_255;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lvtReg_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  lvtReg_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  lvtReg_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  lvtReg_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  lvtReg_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  lvtReg_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  lvtReg_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  lvtReg_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  lvtReg_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  lvtReg_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  lvtReg_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  lvtReg_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  lvtReg_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  lvtReg_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  lvtReg_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  lvtReg_15 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  lvtReg_16 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  lvtReg_17 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  lvtReg_18 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  lvtReg_19 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  lvtReg_20 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  lvtReg_21 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  lvtReg_22 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  lvtReg_23 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  lvtReg_24 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  lvtReg_25 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  lvtReg_26 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  lvtReg_27 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  lvtReg_28 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  lvtReg_29 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  lvtReg_30 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  lvtReg_31 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  lvtReg_32 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  lvtReg_33 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  lvtReg_34 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  lvtReg_35 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  lvtReg_36 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  lvtReg_37 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  lvtReg_38 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  lvtReg_39 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  lvtReg_40 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  lvtReg_41 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  lvtReg_42 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  lvtReg_43 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  lvtReg_44 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  lvtReg_45 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  lvtReg_46 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  lvtReg_47 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  lvtReg_48 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  lvtReg_49 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  lvtReg_50 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  lvtReg_51 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  lvtReg_52 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  lvtReg_53 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  lvtReg_54 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  lvtReg_55 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  lvtReg_56 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  lvtReg_57 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  lvtReg_58 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  lvtReg_59 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  lvtReg_60 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  lvtReg_61 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  lvtReg_62 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  lvtReg_63 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  lvtReg_64 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  lvtReg_65 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  lvtReg_66 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  lvtReg_67 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  lvtReg_68 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  lvtReg_69 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  lvtReg_70 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  lvtReg_71 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  lvtReg_72 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  lvtReg_73 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  lvtReg_74 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  lvtReg_75 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  lvtReg_76 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  lvtReg_77 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  lvtReg_78 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  lvtReg_79 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  lvtReg_80 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  lvtReg_81 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  lvtReg_82 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  lvtReg_83 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  lvtReg_84 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  lvtReg_85 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  lvtReg_86 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  lvtReg_87 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  lvtReg_88 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  lvtReg_89 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  lvtReg_90 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  lvtReg_91 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  lvtReg_92 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  lvtReg_93 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  lvtReg_94 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  lvtReg_95 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  lvtReg_96 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  lvtReg_97 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  lvtReg_98 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  lvtReg_99 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  lvtReg_100 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  lvtReg_101 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  lvtReg_102 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  lvtReg_103 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  lvtReg_104 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  lvtReg_105 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  lvtReg_106 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  lvtReg_107 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  lvtReg_108 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  lvtReg_109 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  lvtReg_110 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  lvtReg_111 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  lvtReg_112 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  lvtReg_113 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  lvtReg_114 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  lvtReg_115 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  lvtReg_116 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  lvtReg_117 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  lvtReg_118 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  lvtReg_119 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  lvtReg_120 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  lvtReg_121 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  lvtReg_122 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  lvtReg_123 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  lvtReg_124 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  lvtReg_125 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  lvtReg_126 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  lvtReg_127 = _RAND_127[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LVTMultiPortRams(
  input        clock,
  input        reset,
  input  [9:0] io_wrAddr_0,
  input  [9:0] io_wrAddr_1,
  input  [7:0] io_wrData_0,
  input  [7:0] io_wrData_1,
  input        io_wrEna_0,
  input        io_wrEna_1,
  input  [9:0] io_rdAddr_0,
  input  [9:0] io_rdAddr_1,
  output [7:0] io_rdData_0,
  output [7:0] io_rdData_1
);
  wire  Memory_clock; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_io_rdAddr; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_io_rdData; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_io_wrEna; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_io_wrData; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_io_wrAddr; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_1_clock; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_1_io_rdAddr; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_1_io_rdData; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_1_io_wrEna; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_1_io_wrData; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_1_io_wrAddr; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_2_clock; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_2_io_rdAddr; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_2_io_rdData; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_2_io_wrEna; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_2_io_wrData; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_2_io_wrAddr; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_3_clock; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_3_io_rdAddr; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_3_io_rdData; // @[LVTMultiPortRams.scala 51:44]
  wire  Memory_3_io_wrEna; // @[LVTMultiPortRams.scala 51:44]
  wire [7:0] Memory_3_io_wrData; // @[LVTMultiPortRams.scala 51:44]
  wire [9:0] Memory_3_io_wrAddr; // @[LVTMultiPortRams.scala 51:44]
  wire  lvt_clock; // @[LVTMultiPortRams.scala 52:19]
  wire  lvt_reset; // @[LVTMultiPortRams.scala 52:19]
  wire [9:0] lvt_io_wrAddr_0; // @[LVTMultiPortRams.scala 52:19]
  wire [9:0] lvt_io_wrAddr_1; // @[LVTMultiPortRams.scala 52:19]
  wire  lvt_io_wrEna_0; // @[LVTMultiPortRams.scala 52:19]
  wire  lvt_io_wrEna_1; // @[LVTMultiPortRams.scala 52:19]
  wire [9:0] lvt_io_rdAddr_0; // @[LVTMultiPortRams.scala 52:19]
  wire [9:0] lvt_io_rdAddr_1; // @[LVTMultiPortRams.scala 52:19]
  wire [1:0] lvt_io_rdIdx_0; // @[LVTMultiPortRams.scala 52:19]
  wire [1:0] lvt_io_rdIdx_1; // @[LVTMultiPortRams.scala 52:19]
  wire [3:0] _io_rdData_0_T = lvt_io_rdIdx_0 * 2'h2; // @[LVTMultiPortRams.scala 71:30]
  wire [4:0] _io_rdData_0_T_1 = {{1'd0}, _io_rdData_0_T}; // @[LVTMultiPortRams.scala 71:36]
  wire [7:0] mems_0_rdData = Memory_io_rdData; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 51:21]
  wire [7:0] mems_1_rdData = Memory_1_io_rdData; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 51:21]
  wire [7:0] _GEN_6 = 2'h1 == _io_rdData_0_T_1[1:0] ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 71:18 LVTMultiPortRams.scala 71:18]
  wire [7:0] mems_2_rdData = Memory_2_io_rdData; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 51:21]
  wire [7:0] _GEN_11 = 2'h2 == _io_rdData_0_T_1[1:0] ? mems_2_rdData : _GEN_6; // @[LVTMultiPortRams.scala 71:18 LVTMultiPortRams.scala 71:18]
  wire [7:0] mems_3_rdData = Memory_3_io_rdData; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 51:21]
  wire [3:0] _io_rdData_1_T = lvt_io_rdIdx_1 * 2'h2; // @[LVTMultiPortRams.scala 71:30]
  wire [3:0] _io_rdData_1_T_2 = _io_rdData_1_T + 4'h1; // @[LVTMultiPortRams.scala 71:36]
  wire [7:0] _GEN_26 = 2'h1 == _io_rdData_1_T_2[1:0] ? mems_1_rdData : mems_0_rdData; // @[LVTMultiPortRams.scala 71:18 LVTMultiPortRams.scala 71:18]
  wire [7:0] _GEN_31 = 2'h2 == _io_rdData_1_T_2[1:0] ? mems_2_rdData : _GEN_26; // @[LVTMultiPortRams.scala 71:18 LVTMultiPortRams.scala 71:18]
  Memory Memory ( // @[LVTMultiPortRams.scala 51:44]
    .clock(Memory_clock),
    .io_rdAddr(Memory_io_rdAddr),
    .io_rdData(Memory_io_rdData),
    .io_wrEna(Memory_io_wrEna),
    .io_wrData(Memory_io_wrData),
    .io_wrAddr(Memory_io_wrAddr)
  );
  Memory Memory_1 ( // @[LVTMultiPortRams.scala 51:44]
    .clock(Memory_1_clock),
    .io_rdAddr(Memory_1_io_rdAddr),
    .io_rdData(Memory_1_io_rdData),
    .io_wrEna(Memory_1_io_wrEna),
    .io_wrData(Memory_1_io_wrData),
    .io_wrAddr(Memory_1_io_wrAddr)
  );
  Memory Memory_2 ( // @[LVTMultiPortRams.scala 51:44]
    .clock(Memory_2_clock),
    .io_rdAddr(Memory_2_io_rdAddr),
    .io_rdData(Memory_2_io_rdData),
    .io_wrEna(Memory_2_io_wrEna),
    .io_wrData(Memory_2_io_wrData),
    .io_wrAddr(Memory_2_io_wrAddr)
  );
  Memory Memory_3 ( // @[LVTMultiPortRams.scala 51:44]
    .clock(Memory_3_clock),
    .io_rdAddr(Memory_3_io_rdAddr),
    .io_rdData(Memory_3_io_rdData),
    .io_wrEna(Memory_3_io_wrEna),
    .io_wrData(Memory_3_io_wrData),
    .io_wrAddr(Memory_3_io_wrAddr)
  );
  LiveValueTable lvt ( // @[LVTMultiPortRams.scala 52:19]
    .clock(lvt_clock),
    .reset(lvt_reset),
    .io_wrAddr_0(lvt_io_wrAddr_0),
    .io_wrAddr_1(lvt_io_wrAddr_1),
    .io_wrEna_0(lvt_io_wrEna_0),
    .io_wrEna_1(lvt_io_wrEna_1),
    .io_rdAddr_0(lvt_io_rdAddr_0),
    .io_rdAddr_1(lvt_io_rdAddr_1),
    .io_rdIdx_0(lvt_io_rdIdx_0),
    .io_rdIdx_1(lvt_io_rdIdx_1)
  );
  assign io_rdData_0 = 2'h3 == _io_rdData_0_T_1[1:0] ? mems_3_rdData : _GEN_11; // @[LVTMultiPortRams.scala 71:18 LVTMultiPortRams.scala 71:18]
  assign io_rdData_1 = 2'h3 == _io_rdData_1_T_2[1:0] ? mems_3_rdData : _GEN_31; // @[LVTMultiPortRams.scala 71:18 LVTMultiPortRams.scala 71:18]
  assign Memory_clock = clock;
  assign Memory_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 59:30]
  assign Memory_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 56:29]
  assign Memory_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 58:30]
  assign Memory_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 57:30]
  assign Memory_1_clock = clock;
  assign Memory_1_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 59:30]
  assign Memory_1_io_wrEna = io_wrEna_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 56:29]
  assign Memory_1_io_wrData = io_wrData_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 58:30]
  assign Memory_1_io_wrAddr = io_wrAddr_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 57:30]
  assign Memory_2_clock = clock;
  assign Memory_2_io_rdAddr = io_rdAddr_0; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 59:30]
  assign Memory_2_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 56:29]
  assign Memory_2_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 58:30]
  assign Memory_2_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 57:30]
  assign Memory_3_clock = clock;
  assign Memory_3_io_rdAddr = io_rdAddr_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 59:30]
  assign Memory_3_io_wrEna = io_wrEna_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 56:29]
  assign Memory_3_io_wrData = io_wrData_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 58:30]
  assign Memory_3_io_wrAddr = io_wrAddr_1; // @[LVTMultiPortRams.scala 51:21 LVTMultiPortRams.scala 57:30]
  assign lvt_clock = clock;
  assign lvt_reset = reset;
  assign lvt_io_wrAddr_0 = io_wrAddr_0; // @[LVTMultiPortRams.scala 64:22]
  assign lvt_io_wrAddr_1 = io_wrAddr_1; // @[LVTMultiPortRams.scala 64:22]
  assign lvt_io_wrEna_0 = io_wrEna_0; // @[LVTMultiPortRams.scala 63:21]
  assign lvt_io_wrEna_1 = io_wrEna_1; // @[LVTMultiPortRams.scala 63:21]
  assign lvt_io_rdAddr_0 = io_rdAddr_0; // @[LVTMultiPortRams.scala 67:22]
  assign lvt_io_rdAddr_1 = io_rdAddr_1; // @[LVTMultiPortRams.scala 67:22]
endmodule
